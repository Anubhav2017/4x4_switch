-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity inputPort_1_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    in_data_1_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_1_pipe_read_data : in   std_logic_vector(31 downto 0);
    noblock_obuf_1_3_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_3_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_1_4_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_4_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_1_1_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_1_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_1_2_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_2_pipe_write_data : out  std_logic_vector(32 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity inputPort_1_Daemon;
architecture inputPort_1_Daemon_arch of inputPort_1_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal inputPort_1_Daemon_CP_3_start: Boolean;
  signal inputPort_1_Daemon_CP_3_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal phi_stmt_67_req_1 : boolean;
  signal do_while_stmt_65_branch_req_0 : boolean;
  signal phi_stmt_76_req_0 : boolean;
  signal phi_stmt_76_ack_0 : boolean;
  signal phi_stmt_67_req_0 : boolean;
  signal phi_stmt_67_ack_0 : boolean;
  signal next_count_down_103_72_buf_req_0 : boolean;
  signal next_count_down_103_72_buf_ack_0 : boolean;
  signal next_count_down_103_72_buf_req_1 : boolean;
  signal next_count_down_103_72_buf_ack_1 : boolean;
  signal RPIPE_in_data_1_75_inst_req_0 : boolean;
  signal RPIPE_in_data_1_75_inst_ack_0 : boolean;
  signal RPIPE_in_data_1_75_inst_req_1 : boolean;
  signal RPIPE_in_data_1_75_inst_ack_1 : boolean;
  signal phi_stmt_76_req_1 : boolean;
  signal next_last_dest_id_109_79_buf_req_0 : boolean;
  signal next_last_dest_id_109_79_buf_ack_0 : boolean;
  signal next_last_dest_id_109_79_buf_req_1 : boolean;
  signal next_last_dest_id_109_79_buf_ack_1 : boolean;
  signal WPIPE_noblock_obuf_1_1_121_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_1_1_121_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_1_1_121_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_1_1_121_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_1_2_130_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_1_2_130_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_1_2_130_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_1_2_130_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_1_3_139_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_1_3_139_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_1_3_139_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_1_3_139_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_1_4_148_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_1_4_148_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_1_4_148_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_1_4_148_inst_ack_1 : boolean;
  signal do_while_stmt_65_branch_ack_0 : boolean;
  signal do_while_stmt_65_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "inputPort_1_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  inputPort_1_Daemon_CP_3_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "inputPort_1_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_1_Daemon_CP_3_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= inputPort_1_Daemon_CP_3_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_1_Daemon_CP_3_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  inputPort_1_Daemon_CP_3: Block -- control-path 
    signal inputPort_1_Daemon_CP_3_elements: BooleanArray(72 downto 0);
    -- 
  begin -- 
    inputPort_1_Daemon_CP_3_elements(0) <= inputPort_1_Daemon_CP_3_start;
    inputPort_1_Daemon_CP_3_symbol <= inputPort_1_Daemon_CP_3_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_64/$entry
      -- CP-element group 0: 	 branch_block_stmt_64/branch_block_stmt_64__entry__
      -- CP-element group 0: 	 branch_block_stmt_64/do_while_stmt_65__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	72 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_64/$exit
      -- CP-element group 1: 	 branch_block_stmt_64/branch_block_stmt_64__exit__
      -- CP-element group 1: 	 branch_block_stmt_64/do_while_stmt_65__exit__
      -- 
    inputPort_1_Daemon_CP_3_elements(1) <= inputPort_1_Daemon_CP_3_elements(72);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_64/do_while_stmt_65/$entry
      -- CP-element group 2: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65__entry__
      -- 
    inputPort_1_Daemon_CP_3_elements(2) <= inputPort_1_Daemon_CP_3_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	72 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65__exit__
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_64/do_while_stmt_65/loop_back
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	71 
    -- CP-element group 5: 	70 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_64/do_while_stmt_65/condition_done
      -- CP-element group 5: 	 branch_block_stmt_64/do_while_stmt_65/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_64/do_while_stmt_65/loop_taken/$entry
      -- 
    inputPort_1_Daemon_CP_3_elements(5) <= inputPort_1_Daemon_CP_3_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	69 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_64/do_while_stmt_65/loop_body_done
      -- 
    inputPort_1_Daemon_CP_3_elements(6) <= inputPort_1_Daemon_CP_3_elements(69);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	43 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/back_edge_to_loop_body
      -- 
    inputPort_1_Daemon_CP_3_elements(7) <= inputPort_1_Daemon_CP_3_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	45 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/first_time_through_loop_body
      -- 
    inputPort_1_Daemon_CP_3_elements(8) <= inputPort_1_Daemon_CP_3_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	68 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	37 
    -- CP-element group 9: 	38 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_73_sample_start_
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	68 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/condition_evaluated
      -- 
    condition_evaluated_27_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_27_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(10), ack => do_while_stmt_65_branch_req_0); -- 
    inputPort_1_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(14) & inputPort_1_Daemon_CP_3_elements(68);
      gj_inputPort_1_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	37 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11: 	39 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_sample_start__ps
      -- 
    inputPort_1_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(9) & inputPort_1_Daemon_CP_3_elements(15) & inputPort_1_Daemon_CP_3_elements(37) & inputPort_1_Daemon_CP_3_elements(14);
      gj_inputPort_1_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	40 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	69 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	37 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_73_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_sample_completed_
      -- 
    inputPort_1_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(17) & inputPort_1_Daemon_CP_3_elements(35) & inputPort_1_Daemon_CP_3_elements(40);
      gj_inputPort_1_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	32 
    -- CP-element group 13: 	38 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13: 	41 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_update_start__ps
      -- 
    inputPort_1_Daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(16) & inputPort_1_Daemon_CP_3_elements(32) & inputPort_1_Daemon_CP_3_elements(38);
      gj_inputPort_1_Daemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	36 
    -- CP-element group 14: 	42 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/aggregated_phi_update_ack
      -- 
    inputPort_1_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(18) & inputPort_1_Daemon_CP_3_elements(36) & inputPort_1_Daemon_CP_3_elements(42);
      gj_inputPort_1_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_sample_start_
      -- 
    inputPort_1_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(9) & inputPort_1_Daemon_CP_3_elements(12);
      gj_inputPort_1_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	57 
    -- CP-element group 16: 	66 
    -- CP-element group 16: 	63 
    -- CP-element group 16: 	60 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_update_start_
      -- 
    inputPort_1_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(9) & inputPort_1_Daemon_CP_3_elements(57) & inputPort_1_Daemon_CP_3_elements(66) & inputPort_1_Daemon_CP_3_elements(63) & inputPort_1_Daemon_CP_3_elements(60);
      gj_inputPort_1_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_sample_completed__ps
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	65 
    -- CP-element group 18: 	56 
    -- CP-element group 18: 	59 
    -- CP-element group 18: 	62 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_update_completed__ps
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_loopback_trigger
      -- 
    inputPort_1_Daemon_CP_3_elements(19) <= inputPort_1_Daemon_CP_3_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_loopback_sample_req_ps
      -- 
    phi_stmt_67_loopback_sample_req_42_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_67_loopback_sample_req_42_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(20), ack => phi_stmt_67_req_1); -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_entry_trigger
      -- 
    inputPort_1_Daemon_CP_3_elements(21) <= inputPort_1_Daemon_CP_3_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_entry_sample_req_ps
      -- 
    phi_stmt_67_entry_sample_req_45_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_67_entry_sample_req_45_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(22), ack => phi_stmt_67_req_0); -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_phi_mux_ack_ps
      -- 
    phi_stmt_67_phi_mux_ack_48_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_67_ack_0, ack => inputPort_1_Daemon_CP_3_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/type_cast_71_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/type_cast_71_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/type_cast_71_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/type_cast_71_sample_completed_
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/type_cast_71_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/type_cast_71_update_start_
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/type_cast_71_update_completed__ps
      -- 
    inputPort_1_Daemon_CP_3_elements(26) <= inputPort_1_Daemon_CP_3_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/type_cast_71_update_completed_
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => inputPort_1_Daemon_CP_3_elements(25), ack => inputPort_1_Daemon_CP_3_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_72_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_72_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_72_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_72_Sample/req
      -- 
    req_69_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_69_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(28), ack => next_count_down_103_72_buf_req_0); -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_72_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_72_update_start_
      -- CP-element group 29: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_72_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_72_Update/req
      -- 
    req_74_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_74_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(29), ack => next_count_down_103_72_buf_req_1); -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_72_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_72_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_72_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_72_Sample/ack
      -- 
    ack_70_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_103_72_buf_ack_0, ack => inputPort_1_Daemon_CP_3_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_72_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_72_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_72_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_72_Update/ack
      -- 
    ack_75_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_103_72_buf_ack_1, ack => inputPort_1_Daemon_CP_3_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	57 
    -- CP-element group 32: 	66 
    -- CP-element group 32: 	63 
    -- CP-element group 32: 	60 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_73_update_start_
      -- 
    inputPort_1_Daemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(9) & inputPort_1_Daemon_CP_3_elements(57) & inputPort_1_Daemon_CP_3_elements(66) & inputPort_1_Daemon_CP_3_elements(63) & inputPort_1_Daemon_CP_3_elements(60);
      gj_inputPort_1_Daemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/RPIPE_in_data_1_75_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/RPIPE_in_data_1_75_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/RPIPE_in_data_1_75_Sample/rr
      -- 
    rr_88_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_88_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(33), ack => RPIPE_in_data_1_75_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(11) & inputPort_1_Daemon_CP_3_elements(36);
      gj_inputPort_1_Daemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	13 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/RPIPE_in_data_1_75_update_start_
      -- CP-element group 34: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/RPIPE_in_data_1_75_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/RPIPE_in_data_1_75_Update/cr
      -- 
    cr_93_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_93_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(34), ack => RPIPE_in_data_1_75_inst_req_1); -- 
    inputPort_1_Daemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(13) & inputPort_1_Daemon_CP_3_elements(35);
      gj_inputPort_1_Daemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/RPIPE_in_data_1_75_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/RPIPE_in_data_1_75_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/RPIPE_in_data_1_75_Sample/ra
      -- 
    ra_89_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_1_75_inst_ack_0, ack => inputPort_1_Daemon_CP_3_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	65 
    -- CP-element group 36: 	56 
    -- CP-element group 36: 	59 
    -- CP-element group 36: 	62 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_73_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/RPIPE_in_data_1_75_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/RPIPE_in_data_1_75_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/RPIPE_in_data_1_75_Update/ca
      -- 
    ca_94_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_1_75_inst_ack_1, ack => inputPort_1_Daemon_CP_3_elements(36)); -- 
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	9 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	12 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	11 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_sample_start_
      -- 
    inputPort_1_Daemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(9) & inputPort_1_Daemon_CP_3_elements(12);
      gj_inputPort_1_Daemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	9 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	57 
    -- CP-element group 38: 	66 
    -- CP-element group 38: 	63 
    -- CP-element group 38: 	60 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	13 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_update_start_
      -- 
    inputPort_1_Daemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(9) & inputPort_1_Daemon_CP_3_elements(57) & inputPort_1_Daemon_CP_3_elements(66) & inputPort_1_Daemon_CP_3_elements(63) & inputPort_1_Daemon_CP_3_elements(60);
      gj_inputPort_1_Daemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	11 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_sample_start__ps
      -- 
    inputPort_1_Daemon_CP_3_elements(39) <= inputPort_1_Daemon_CP_3_elements(11);
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	12 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_sample_completed__ps
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	13 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_update_start__ps
      -- 
    inputPort_1_Daemon_CP_3_elements(41) <= inputPort_1_Daemon_CP_3_elements(13);
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	14 
    -- CP-element group 42: 	65 
    -- CP-element group 42: 	56 
    -- CP-element group 42: 	59 
    -- CP-element group 42: 	62 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_update_completed__ps
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	7 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_loopback_trigger
      -- 
    inputPort_1_Daemon_CP_3_elements(43) <= inputPort_1_Daemon_CP_3_elements(7);
    -- CP-element group 44:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_loopback_sample_req
      -- CP-element group 44: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_loopback_sample_req_ps
      -- 
    phi_stmt_76_loopback_sample_req_104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_76_loopback_sample_req_104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(44), ack => phi_stmt_76_req_1); -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	8 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_entry_trigger
      -- 
    inputPort_1_Daemon_CP_3_elements(45) <= inputPort_1_Daemon_CP_3_elements(8);
    -- CP-element group 46:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_entry_sample_req
      -- CP-element group 46: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_entry_sample_req_ps
      -- 
    phi_stmt_76_entry_sample_req_107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_76_entry_sample_req_107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(46), ack => phi_stmt_76_req_0); -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_phi_mux_ack
      -- CP-element group 47: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_phi_mux_ack_ps
      -- 
    phi_stmt_76_phi_mux_ack_110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_76_ack_0, ack => inputPort_1_Daemon_CP_3_elements(47)); -- 
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/konst_78_sample_start__ps
      -- CP-element group 48: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/konst_78_sample_completed__ps
      -- CP-element group 48: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/konst_78_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/konst_78_sample_completed_
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/konst_78_update_start__ps
      -- CP-element group 49: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/konst_78_update_start_
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/konst_78_update_completed__ps
      -- 
    inputPort_1_Daemon_CP_3_elements(50) <= inputPort_1_Daemon_CP_3_elements(51);
    -- CP-element group 51:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	50 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/konst_78_update_completed_
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(51) is a control-delay.
    cp_element_51_delay: control_delay_element  generic map(name => " 51_delay", delay_value => 1)  port map(req => inputPort_1_Daemon_CP_3_elements(49), ack => inputPort_1_Daemon_CP_3_elements(51), clk => clk, reset =>reset);
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_Sample/req
      -- 
    req_131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(52), ack => next_last_dest_id_109_79_buf_req_0); -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_update_start_
      -- CP-element group 53: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_Update/req
      -- 
    req_136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(53), ack => next_last_dest_id_109_79_buf_req_1); -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_Sample/ack
      -- 
    ack_132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_109_79_buf_ack_0, ack => inputPort_1_Daemon_CP_3_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_Update/ack
      -- 
    ack_137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_109_79_buf_ack_1, ack => inputPort_1_Daemon_CP_3_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	18 
    -- CP-element group 56: 	36 
    -- CP-element group 56: 	42 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_1_121_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_1_121_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_1_121_Sample/req
      -- 
    req_146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(56), ack => WPIPE_noblock_obuf_1_1_121_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(18) & inputPort_1_Daemon_CP_3_elements(36) & inputPort_1_Daemon_CP_3_elements(42) & inputPort_1_Daemon_CP_3_elements(58);
      gj_inputPort_1_Daemon_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	16 
    -- CP-element group 57: 	32 
    -- CP-element group 57: 	38 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_1_121_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_1_121_update_start_
      -- CP-element group 57: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_1_121_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_1_121_Sample/ack
      -- CP-element group 57: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_1_121_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_1_121_Update/req
      -- 
    ack_147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_1_121_inst_ack_0, ack => inputPort_1_Daemon_CP_3_elements(57)); -- 
    req_151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(57), ack => WPIPE_noblock_obuf_1_1_121_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	69 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_1_121_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_1_121_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_1_121_Update/ack
      -- 
    ack_152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_1_121_inst_ack_1, ack => inputPort_1_Daemon_CP_3_elements(58)); -- 
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	18 
    -- CP-element group 59: 	36 
    -- CP-element group 59: 	42 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_2_130_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_2_130_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_2_130_Sample/req
      -- 
    req_160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(59), ack => WPIPE_noblock_obuf_1_2_130_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(18) & inputPort_1_Daemon_CP_3_elements(36) & inputPort_1_Daemon_CP_3_elements(42) & inputPort_1_Daemon_CP_3_elements(61);
      gj_inputPort_1_Daemon_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	16 
    -- CP-element group 60: 	32 
    -- CP-element group 60: 	38 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_2_130_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_2_130_update_start_
      -- CP-element group 60: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_2_130_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_2_130_Sample/ack
      -- CP-element group 60: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_2_130_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_2_130_Update/req
      -- 
    ack_161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_2_130_inst_ack_0, ack => inputPort_1_Daemon_CP_3_elements(60)); -- 
    req_165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(60), ack => WPIPE_noblock_obuf_1_2_130_inst_req_1); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	69 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_2_130_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_2_130_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_2_130_Update/ack
      -- 
    ack_166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_2_130_inst_ack_1, ack => inputPort_1_Daemon_CP_3_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	18 
    -- CP-element group 62: 	36 
    -- CP-element group 62: 	42 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_3_139_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_3_139_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_3_139_Sample/req
      -- 
    req_174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(62), ack => WPIPE_noblock_obuf_1_3_139_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(18) & inputPort_1_Daemon_CP_3_elements(36) & inputPort_1_Daemon_CP_3_elements(42) & inputPort_1_Daemon_CP_3_elements(64);
      gj_inputPort_1_Daemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	16 
    -- CP-element group 63: 	32 
    -- CP-element group 63: 	38 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_3_139_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_3_139_update_start_
      -- CP-element group 63: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_3_139_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_3_139_Sample/ack
      -- CP-element group 63: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_3_139_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_3_139_Update/req
      -- 
    ack_175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_3_139_inst_ack_0, ack => inputPort_1_Daemon_CP_3_elements(63)); -- 
    req_179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(63), ack => WPIPE_noblock_obuf_1_3_139_inst_req_1); -- 
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	69 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_3_139_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_3_139_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_3_139_Update/ack
      -- 
    ack_180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_3_139_inst_ack_1, ack => inputPort_1_Daemon_CP_3_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	18 
    -- CP-element group 65: 	36 
    -- CP-element group 65: 	42 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_4_148_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_4_148_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_4_148_Sample/req
      -- 
    req_188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(65), ack => WPIPE_noblock_obuf_1_4_148_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(18) & inputPort_1_Daemon_CP_3_elements(36) & inputPort_1_Daemon_CP_3_elements(42) & inputPort_1_Daemon_CP_3_elements(67);
      gj_inputPort_1_Daemon_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	16 
    -- CP-element group 66: 	32 
    -- CP-element group 66: 	38 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_4_148_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_4_148_update_start_
      -- CP-element group 66: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_4_148_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_4_148_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_4_148_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_4_148_Update/req
      -- 
    ack_189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_4_148_inst_ack_0, ack => inputPort_1_Daemon_CP_3_elements(66)); -- 
    req_193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(66), ack => WPIPE_noblock_obuf_1_4_148_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_4_148_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_4_148_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_4_148_Update/ack
      -- 
    ack_194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_4_148_inst_ack_1, ack => inputPort_1_Daemon_CP_3_elements(67)); -- 
    -- CP-element group 68:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	9 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	10 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(68) is a control-delay.
    cp_element_68_delay: control_delay_element  generic map(name => " 68_delay", delay_value => 1)  port map(req => inputPort_1_Daemon_CP_3_elements(9), ack => inputPort_1_Daemon_CP_3_elements(68), clk => clk, reset =>reset);
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	12 
    -- CP-element group 69: 	61 
    -- CP-element group 69: 	58 
    -- CP-element group 69: 	64 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	6 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/$exit
      -- 
    inputPort_1_Daemon_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(12) & inputPort_1_Daemon_CP_3_elements(61) & inputPort_1_Daemon_CP_3_elements(58) & inputPort_1_Daemon_CP_3_elements(64) & inputPort_1_Daemon_CP_3_elements(67);
      gj_inputPort_1_Daemon_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	5 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_64/do_while_stmt_65/loop_exit/$exit
      -- CP-element group 70: 	 branch_block_stmt_64/do_while_stmt_65/loop_exit/ack
      -- 
    ack_199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_65_branch_ack_0, ack => inputPort_1_Daemon_CP_3_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	5 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_64/do_while_stmt_65/loop_taken/$exit
      -- CP-element group 71: 	 branch_block_stmt_64/do_while_stmt_65/loop_taken/ack
      -- 
    ack_203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_65_branch_ack_1, ack => inputPort_1_Daemon_CP_3_elements(71)); -- 
    -- CP-element group 72:  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	3 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	1 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_64/do_while_stmt_65/$exit
      -- 
    inputPort_1_Daemon_CP_3_elements(72) <= inputPort_1_Daemon_CP_3_elements(3);
    inputPort_1_Daemon_do_while_stmt_65_terminator_204: loop_terminator -- 
      generic map (name => " inputPort_1_Daemon_do_while_stmt_65_terminator_204", max_iterations_in_flight =>7) 
      port map(loop_body_exit => inputPort_1_Daemon_CP_3_elements(6),loop_continue => inputPort_1_Daemon_CP_3_elements(71),loop_terminate => inputPort_1_Daemon_CP_3_elements(70),loop_back => inputPort_1_Daemon_CP_3_elements(4),loop_exit => inputPort_1_Daemon_CP_3_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_67_phi_seq_76_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_1_Daemon_CP_3_elements(21);
      inputPort_1_Daemon_CP_3_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_1_Daemon_CP_3_elements(24);
      inputPort_1_Daemon_CP_3_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_1_Daemon_CP_3_elements(26);
      inputPort_1_Daemon_CP_3_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_1_Daemon_CP_3_elements(19);
      inputPort_1_Daemon_CP_3_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_1_Daemon_CP_3_elements(30);
      inputPort_1_Daemon_CP_3_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_1_Daemon_CP_3_elements(31);
      inputPort_1_Daemon_CP_3_elements(20) <= phi_mux_reqs(1);
      phi_stmt_67_phi_seq_76 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_67_phi_seq_76") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_1_Daemon_CP_3_elements(11), 
          phi_sample_ack => inputPort_1_Daemon_CP_3_elements(17), 
          phi_update_req => inputPort_1_Daemon_CP_3_elements(13), 
          phi_update_ack => inputPort_1_Daemon_CP_3_elements(18), 
          phi_mux_ack => inputPort_1_Daemon_CP_3_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_76_phi_seq_138_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_1_Daemon_CP_3_elements(45);
      inputPort_1_Daemon_CP_3_elements(48)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_1_Daemon_CP_3_elements(48);
      inputPort_1_Daemon_CP_3_elements(49)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_1_Daemon_CP_3_elements(50);
      inputPort_1_Daemon_CP_3_elements(46) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_1_Daemon_CP_3_elements(43);
      inputPort_1_Daemon_CP_3_elements(52)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_1_Daemon_CP_3_elements(54);
      inputPort_1_Daemon_CP_3_elements(53)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_1_Daemon_CP_3_elements(55);
      inputPort_1_Daemon_CP_3_elements(44) <= phi_mux_reqs(1);
      phi_stmt_76_phi_seq_138 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_76_phi_seq_138") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_1_Daemon_CP_3_elements(39), 
          phi_sample_ack => inputPort_1_Daemon_CP_3_elements(40), 
          phi_update_req => inputPort_1_Daemon_CP_3_elements(41), 
          phi_update_ack => inputPort_1_Daemon_CP_3_elements(42), 
          phi_mux_ack => inputPort_1_Daemon_CP_3_elements(47), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_28_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= inputPort_1_Daemon_CP_3_elements(7);
        preds(1)  <= inputPort_1_Daemon_CP_3_elements(8);
        entry_tmerge_28 : transition_merge -- 
          generic map(name => " entry_tmerge_28")
          port map (preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal RPIPE_in_data_1_75_wire : std_logic_vector(31 downto 0);
    signal R_ONE_1_111_wire_constant : std_logic_vector(0 downto 0);
    signal SUB_u16_u16_101_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_98_wire : std_logic_vector(15 downto 0);
    signal count_down_67 : std_logic_vector(15 downto 0);
    signal data_to_outport_114 : std_logic_vector(32 downto 0);
    signal dest_id_89 : std_logic_vector(7 downto 0);
    signal input_word_73 : std_logic_vector(31 downto 0);
    signal konst_100_wire_constant : std_logic_vector(15 downto 0);
    signal konst_117_wire_constant : std_logic_vector(7 downto 0);
    signal konst_126_wire_constant : std_logic_vector(7 downto 0);
    signal konst_135_wire_constant : std_logic_vector(7 downto 0);
    signal konst_144_wire_constant : std_logic_vector(7 downto 0);
    signal konst_152_wire_constant : std_logic_vector(0 downto 0);
    signal konst_78_wire_constant : std_logic_vector(7 downto 0);
    signal konst_83_wire_constant : std_logic_vector(15 downto 0);
    signal konst_97_wire_constant : std_logic_vector(15 downto 0);
    signal last_dest_id_76 : std_logic_vector(7 downto 0);
    signal new_packet_85 : std_logic_vector(0 downto 0);
    signal next_count_down_103 : std_logic_vector(15 downto 0);
    signal next_count_down_103_72_buffered : std_logic_vector(15 downto 0);
    signal next_last_dest_id_109 : std_logic_vector(7 downto 0);
    signal next_last_dest_id_109_79_buffered : std_logic_vector(7 downto 0);
    signal pkt_length_93 : std_logic_vector(15 downto 0);
    signal send_to_1_119 : std_logic_vector(0 downto 0);
    signal send_to_2_128 : std_logic_vector(0 downto 0);
    signal send_to_3_137 : std_logic_vector(0 downto 0);
    signal send_to_4_146 : std_logic_vector(0 downto 0);
    signal type_cast_71_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    R_ONE_1_111_wire_constant <= "1";
    konst_100_wire_constant <= "0000000000000001";
    konst_117_wire_constant <= "00000001";
    konst_126_wire_constant <= "00000010";
    konst_135_wire_constant <= "00000011";
    konst_144_wire_constant <= "00000100";
    konst_152_wire_constant <= "1";
    konst_78_wire_constant <= "00000000";
    konst_83_wire_constant <= "0000000000000000";
    konst_97_wire_constant <= "0000000000000001";
    type_cast_71_wire_constant <= "0000000000000000";
    phi_stmt_67: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_71_wire_constant & next_count_down_103_72_buffered;
      req <= phi_stmt_67_req_0 & phi_stmt_67_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_67",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_67_ack_0,
          idata => idata,
          odata => count_down_67,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_67
    phi_stmt_76: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_78_wire_constant & next_last_dest_id_109_79_buffered;
      req <= phi_stmt_76_req_0 & phi_stmt_76_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_76",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_76_ack_0,
          idata => idata,
          odata => last_dest_id_76,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_76
    -- flow-through select operator MUX_102_inst
    next_count_down_103 <= SUB_u16_u16_98_wire when (new_packet_85(0) /=  '0') else SUB_u16_u16_101_wire;
    -- flow-through select operator MUX_108_inst
    next_last_dest_id_109 <= dest_id_89 when (new_packet_85(0) /=  '0') else last_dest_id_76;
    -- flow-through slice operator slice_88_inst
    dest_id_89 <= input_word_73(31 downto 24);
    -- flow-through slice operator slice_92_inst
    pkt_length_93 <= input_word_73(23 downto 8);
    next_count_down_103_72_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_count_down_103_72_buf_req_0;
      next_count_down_103_72_buf_ack_0<= wack(0);
      rreq(0) <= next_count_down_103_72_buf_req_1;
      next_count_down_103_72_buf_ack_1<= rack(0);
      next_count_down_103_72_buf : InterlockBuffer generic map ( -- 
        name => "next_count_down_103_72_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_count_down_103,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_count_down_103_72_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_last_dest_id_109_79_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_last_dest_id_109_79_buf_req_0;
      next_last_dest_id_109_79_buf_ack_0<= wack(0);
      rreq(0) <= next_last_dest_id_109_79_buf_req_1;
      next_last_dest_id_109_79_buf_ack_1<= rack(0);
      next_last_dest_id_109_79_buf : InterlockBuffer generic map ( -- 
        name => "next_last_dest_id_109_79_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_last_dest_id_109,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_last_dest_id_109_79_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_73
    process(RPIPE_in_data_1_75_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := RPIPE_in_data_1_75_wire(31 downto 0);
      input_word_73 <= tmp_var; -- 
    end process;
    do_while_stmt_65_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_152_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_65_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_65_branch_req_0,
          ack0 => do_while_stmt_65_branch_ack_0,
          ack1 => do_while_stmt_65_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator CONCAT_u1_u33_113_inst
    process(R_ONE_1_111_wire_constant, input_word_73) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ONE_1_111_wire_constant, input_word_73, tmp_var);
      data_to_outport_114 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_84_inst
    process(count_down_67) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(count_down_67, konst_83_wire_constant, tmp_var);
      new_packet_85 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_118_inst
    process(next_last_dest_id_109) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_109, konst_117_wire_constant, tmp_var);
      send_to_1_119 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_127_inst
    process(next_last_dest_id_109) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_109, konst_126_wire_constant, tmp_var);
      send_to_2_128 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_136_inst
    process(next_last_dest_id_109) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_109, konst_135_wire_constant, tmp_var);
      send_to_3_137 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_145_inst
    process(next_last_dest_id_109) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_109, konst_144_wire_constant, tmp_var);
      send_to_4_146 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_101_inst
    process(count_down_67) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(count_down_67, konst_100_wire_constant, tmp_var);
      SUB_u16_u16_101_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_98_inst
    process(pkt_length_93) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(pkt_length_93, konst_97_wire_constant, tmp_var);
      SUB_u16_u16_98_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_in_data_1_75_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_in_data_1_75_inst_req_0;
      RPIPE_in_data_1_75_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_in_data_1_75_inst_req_1;
      RPIPE_in_data_1_75_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_in_data_1_75_wire <= data_out(31 downto 0);
      in_data_1_read_0_gI: SplitGuardInterface generic map(name => "in_data_1_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      in_data_1_read_0: InputPortRevised -- 
        generic map ( name => "in_data_1_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => in_data_1_pipe_read_req(0),
          oack => in_data_1_pipe_read_ack(0),
          odata => in_data_1_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_noblock_obuf_1_1_121_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_1_1_121_inst_req_0;
      WPIPE_noblock_obuf_1_1_121_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_1_1_121_inst_req_1;
      WPIPE_noblock_obuf_1_1_121_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_1_119(0);
      data_in <= data_to_outport_114;
      noblock_obuf_1_1_write_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_1_write_0: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_1_1", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_1_1_pipe_write_req(0),
          oack => noblock_obuf_1_1_pipe_write_ack(0),
          odata => noblock_obuf_1_1_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_noblock_obuf_1_2_130_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_1_2_130_inst_req_0;
      WPIPE_noblock_obuf_1_2_130_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_1_2_130_inst_req_1;
      WPIPE_noblock_obuf_1_2_130_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_2_128(0);
      data_in <= data_to_outport_114;
      noblock_obuf_1_2_write_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_2_write_1: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_1_2", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_1_2_pipe_write_req(0),
          oack => noblock_obuf_1_2_pipe_write_ack(0),
          odata => noblock_obuf_1_2_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_noblock_obuf_1_3_139_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_1_3_139_inst_req_0;
      WPIPE_noblock_obuf_1_3_139_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_1_3_139_inst_req_1;
      WPIPE_noblock_obuf_1_3_139_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_3_137(0);
      data_in <= data_to_outport_114;
      noblock_obuf_1_3_write_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_3_write_2: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_1_3", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_1_3_pipe_write_req(0),
          oack => noblock_obuf_1_3_pipe_write_ack(0),
          odata => noblock_obuf_1_3_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_noblock_obuf_1_4_148_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_1_4_148_inst_req_0;
      WPIPE_noblock_obuf_1_4_148_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_1_4_148_inst_req_1;
      WPIPE_noblock_obuf_1_4_148_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_4_146(0);
      data_in <= data_to_outport_114;
      noblock_obuf_1_4_write_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_4_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_4_write_3: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_1_4", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_1_4_pipe_write_req(0),
          oack => noblock_obuf_1_4_pipe_write_ack(0),
          odata => noblock_obuf_1_4_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end inputPort_1_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity inputPort_2_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    in_data_2_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_2_pipe_read_data : in   std_logic_vector(31 downto 0);
    noblock_obuf_2_1_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_1_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_2_2_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_2_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_2_3_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_3_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_2_4_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_4_pipe_write_data : out  std_logic_vector(32 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity inputPort_2_Daemon;
architecture inputPort_2_Daemon_arch of inputPort_2_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal inputPort_2_Daemon_CP_205_start: Boolean;
  signal inputPort_2_Daemon_CP_205_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_noblock_obuf_2_3_230_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_2_3_230_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_2_3_230_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_2_3_230_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_2_4_239_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_2_4_239_inst_ack_0 : boolean;
  signal do_while_stmt_157_branch_req_0 : boolean;
  signal phi_stmt_159_req_0 : boolean;
  signal phi_stmt_159_req_1 : boolean;
  signal phi_stmt_159_ack_0 : boolean;
  signal next_count_down_194_161_buf_req_0 : boolean;
  signal next_count_down_194_161_buf_ack_0 : boolean;
  signal next_count_down_194_161_buf_req_1 : boolean;
  signal next_count_down_194_161_buf_ack_1 : boolean;
  signal RPIPE_in_data_2_166_inst_req_0 : boolean;
  signal RPIPE_in_data_2_166_inst_ack_0 : boolean;
  signal RPIPE_in_data_2_166_inst_req_1 : boolean;
  signal RPIPE_in_data_2_166_inst_ack_1 : boolean;
  signal phi_stmt_167_req_1 : boolean;
  signal phi_stmt_167_req_0 : boolean;
  signal phi_stmt_167_ack_0 : boolean;
  signal next_last_dest_id_200_170_buf_req_0 : boolean;
  signal next_last_dest_id_200_170_buf_ack_0 : boolean;
  signal next_last_dest_id_200_170_buf_req_1 : boolean;
  signal next_last_dest_id_200_170_buf_ack_1 : boolean;
  signal WPIPE_noblock_obuf_2_1_212_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_2_1_212_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_2_1_212_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_2_1_212_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_2_2_221_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_2_2_221_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_2_2_221_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_2_2_221_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_2_4_239_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_2_4_239_inst_ack_1 : boolean;
  signal do_while_stmt_157_branch_ack_0 : boolean;
  signal do_while_stmt_157_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "inputPort_2_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  inputPort_2_Daemon_CP_205_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "inputPort_2_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_2_Daemon_CP_205_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= inputPort_2_Daemon_CP_205_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_2_Daemon_CP_205_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  inputPort_2_Daemon_CP_205: Block -- control-path 
    signal inputPort_2_Daemon_CP_205_elements: BooleanArray(72 downto 0);
    -- 
  begin -- 
    inputPort_2_Daemon_CP_205_elements(0) <= inputPort_2_Daemon_CP_205_start;
    inputPort_2_Daemon_CP_205_symbol <= inputPort_2_Daemon_CP_205_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_156/$entry
      -- CP-element group 0: 	 branch_block_stmt_156/branch_block_stmt_156__entry__
      -- CP-element group 0: 	 branch_block_stmt_156/do_while_stmt_157__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	72 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_156/$exit
      -- CP-element group 1: 	 branch_block_stmt_156/branch_block_stmt_156__exit__
      -- CP-element group 1: 	 branch_block_stmt_156/do_while_stmt_157__exit__
      -- 
    inputPort_2_Daemon_CP_205_elements(1) <= inputPort_2_Daemon_CP_205_elements(72);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_156/do_while_stmt_157/$entry
      -- CP-element group 2: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157__entry__
      -- 
    inputPort_2_Daemon_CP_205_elements(2) <= inputPort_2_Daemon_CP_205_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	72 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157__exit__
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_156/do_while_stmt_157/loop_back
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	70 
    -- CP-element group 5: 	71 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_156/do_while_stmt_157/condition_done
      -- CP-element group 5: 	 branch_block_stmt_156/do_while_stmt_157/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_156/do_while_stmt_157/loop_taken/$entry
      -- 
    inputPort_2_Daemon_CP_205_elements(5) <= inputPort_2_Daemon_CP_205_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	69 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_156/do_while_stmt_157/loop_body_done
      -- 
    inputPort_2_Daemon_CP_205_elements(6) <= inputPort_2_Daemon_CP_205_elements(69);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	43 
    -- CP-element group 7: 	21 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/back_edge_to_loop_body
      -- 
    inputPort_2_Daemon_CP_205_elements(7) <= inputPort_2_Daemon_CP_205_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	45 
    -- CP-element group 8: 	23 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/first_time_through_loop_body
      -- 
    inputPort_2_Daemon_CP_205_elements(8) <= inputPort_2_Daemon_CP_205_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	68 
    -- CP-element group 9: 	40 
    -- CP-element group 9: 	39 
    -- CP-element group 9: 	34 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_164_sample_start_
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	68 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/condition_evaluated
      -- 
    condition_evaluated_229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(10), ack => do_while_stmt_157_branch_req_0); -- 
    inputPort_2_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(68) & inputPort_2_Daemon_CP_205_elements(14);
      gj_inputPort_2_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	39 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	35 
    -- CP-element group 11: 	17 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_sample_start__ps
      -- 
    inputPort_2_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 7,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(39) & inputPort_2_Daemon_CP_205_elements(9) & inputPort_2_Daemon_CP_205_elements(15) & inputPort_2_Daemon_CP_205_elements(14);
      gj_inputPort_2_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	37 
    -- CP-element group 12: 	41 
    -- CP-element group 12: 	18 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	69 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	39 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_164_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_sample_completed_
      -- 
    inputPort_2_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(37) & inputPort_2_Daemon_CP_205_elements(41) & inputPort_2_Daemon_CP_205_elements(18);
      gj_inputPort_2_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	40 
    -- CP-element group 13: 	34 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	36 
    -- CP-element group 13: 	19 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_update_start__ps
      -- 
    inputPort_2_Daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(40) & inputPort_2_Daemon_CP_205_elements(34) & inputPort_2_Daemon_CP_205_elements(16);
      gj_inputPort_2_Daemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	42 
    -- CP-element group 14: 	38 
    -- CP-element group 14: 	20 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/aggregated_phi_update_ack
      -- 
    inputPort_2_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(42) & inputPort_2_Daemon_CP_205_elements(38) & inputPort_2_Daemon_CP_205_elements(20);
      gj_inputPort_2_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_sample_start_
      -- 
    inputPort_2_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(9) & inputPort_2_Daemon_CP_205_elements(12);
      gj_inputPort_2_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	63 
    -- CP-element group 16: 	57 
    -- CP-element group 16: 	60 
    -- CP-element group 16: 	66 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_update_start_
      -- 
    inputPort_2_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(9) & inputPort_2_Daemon_CP_205_elements(63) & inputPort_2_Daemon_CP_205_elements(57) & inputPort_2_Daemon_CP_205_elements(60) & inputPort_2_Daemon_CP_205_elements(66);
      gj_inputPort_2_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_sample_start__ps
      -- 
    inputPort_2_Daemon_CP_205_elements(17) <= inputPort_2_Daemon_CP_205_elements(11);
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_sample_completed__ps
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_update_start__ps
      -- 
    inputPort_2_Daemon_CP_205_elements(19) <= inputPort_2_Daemon_CP_205_elements(13);
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	56 
    -- CP-element group 20: 	62 
    -- CP-element group 20: 	59 
    -- CP-element group 20: 	65 
    -- CP-element group 20: 	14 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_update_completed__ps
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_loopback_trigger
      -- 
    inputPort_2_Daemon_CP_205_elements(21) <= inputPort_2_Daemon_CP_205_elements(7);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_loopback_sample_req_ps
      -- 
    phi_stmt_159_loopback_sample_req_244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_159_loopback_sample_req_244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(22), ack => phi_stmt_159_req_0); -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_entry_trigger
      -- 
    inputPort_2_Daemon_CP_205_elements(23) <= inputPort_2_Daemon_CP_205_elements(8);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_entry_sample_req
      -- CP-element group 24: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_entry_sample_req_ps
      -- 
    phi_stmt_159_entry_sample_req_247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_159_entry_sample_req_247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(24), ack => phi_stmt_159_req_1); -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_phi_mux_ack_ps
      -- 
    phi_stmt_159_phi_mux_ack_250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_159_ack_0, ack => inputPort_2_Daemon_CP_205_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_sample_start__ps
      -- CP-element group 26: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_Sample/req
      -- 
    req_263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(26), ack => next_count_down_194_161_buf_req_0); -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_update_start_
      -- CP-element group 27: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_Update/req
      -- 
    req_268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(27), ack => next_count_down_194_161_buf_req_1); -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_Sample/ack
      -- 
    ack_264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_194_161_buf_ack_0, ack => inputPort_2_Daemon_CP_205_elements(28)); -- 
    -- CP-element group 29:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_update_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_Update/ack
      -- 
    ack_269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_194_161_buf_ack_1, ack => inputPort_2_Daemon_CP_205_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/type_cast_163_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/type_cast_163_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/type_cast_163_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/type_cast_163_sample_completed_
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/type_cast_163_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/type_cast_163_update_start_
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	33 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/type_cast_163_update_completed__ps
      -- 
    inputPort_2_Daemon_CP_205_elements(32) <= inputPort_2_Daemon_CP_205_elements(33);
    -- CP-element group 33:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	32 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/type_cast_163_update_completed_
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(33) is a control-delay.
    cp_element_33_delay: control_delay_element  generic map(name => " 33_delay", delay_value => 1)  port map(req => inputPort_2_Daemon_CP_205_elements(31), ack => inputPort_2_Daemon_CP_205_elements(33), clk => clk, reset =>reset);
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	9 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	63 
    -- CP-element group 34: 	57 
    -- CP-element group 34: 	60 
    -- CP-element group 34: 	66 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	13 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_164_update_start_
      -- 
    inputPort_2_Daemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(9) & inputPort_2_Daemon_CP_205_elements(63) & inputPort_2_Daemon_CP_205_elements(57) & inputPort_2_Daemon_CP_205_elements(60) & inputPort_2_Daemon_CP_205_elements(66);
      gj_inputPort_2_Daemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	11 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	38 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/RPIPE_in_data_2_166_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/RPIPE_in_data_2_166_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/RPIPE_in_data_2_166_Sample/rr
      -- 
    rr_290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(35), ack => RPIPE_in_data_2_166_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(11) & inputPort_2_Daemon_CP_205_elements(38);
      gj_inputPort_2_Daemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: 	13 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/RPIPE_in_data_2_166_update_start_
      -- CP-element group 36: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/RPIPE_in_data_2_166_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/RPIPE_in_data_2_166_Update/cr
      -- 
    cr_295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(36), ack => RPIPE_in_data_2_166_inst_req_1); -- 
    inputPort_2_Daemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(37) & inputPort_2_Daemon_CP_205_elements(13);
      gj_inputPort_2_Daemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: 	12 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/RPIPE_in_data_2_166_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/RPIPE_in_data_2_166_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/RPIPE_in_data_2_166_Sample/ra
      -- 
    ra_291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_2_166_inst_ack_0, ack => inputPort_2_Daemon_CP_205_elements(37)); -- 
    -- CP-element group 38:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	56 
    -- CP-element group 38: 	62 
    -- CP-element group 38: 	59 
    -- CP-element group 38: 	65 
    -- CP-element group 38: 	14 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	35 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_164_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/RPIPE_in_data_2_166_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/RPIPE_in_data_2_166_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/RPIPE_in_data_2_166_Update/ca
      -- 
    ca_296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_2_166_inst_ack_1, ack => inputPort_2_Daemon_CP_205_elements(38)); -- 
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	9 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	12 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	11 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_sample_start_
      -- 
    inputPort_2_Daemon_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(9) & inputPort_2_Daemon_CP_205_elements(12);
      gj_inputPort_2_Daemon_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	9 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	63 
    -- CP-element group 40: 	57 
    -- CP-element group 40: 	60 
    -- CP-element group 40: 	66 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	13 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_update_start_
      -- 
    inputPort_2_Daemon_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(9) & inputPort_2_Daemon_CP_205_elements(63) & inputPort_2_Daemon_CP_205_elements(57) & inputPort_2_Daemon_CP_205_elements(60) & inputPort_2_Daemon_CP_205_elements(66);
      gj_inputPort_2_Daemon_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	12 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_sample_completed__ps
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	56 
    -- CP-element group 42: 	62 
    -- CP-element group 42: 	59 
    -- CP-element group 42: 	65 
    -- CP-element group 42: 	14 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_update_completed__ps
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	7 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_loopback_trigger
      -- 
    inputPort_2_Daemon_CP_205_elements(43) <= inputPort_2_Daemon_CP_205_elements(7);
    -- CP-element group 44:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_loopback_sample_req
      -- CP-element group 44: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_loopback_sample_req_ps
      -- 
    phi_stmt_167_loopback_sample_req_306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_167_loopback_sample_req_306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(44), ack => phi_stmt_167_req_1); -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	8 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_entry_trigger
      -- 
    inputPort_2_Daemon_CP_205_elements(45) <= inputPort_2_Daemon_CP_205_elements(8);
    -- CP-element group 46:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_entry_sample_req
      -- CP-element group 46: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_entry_sample_req_ps
      -- 
    phi_stmt_167_entry_sample_req_309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_167_entry_sample_req_309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(46), ack => phi_stmt_167_req_0); -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_phi_mux_ack
      -- CP-element group 47: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_phi_mux_ack_ps
      -- 
    phi_stmt_167_phi_mux_ack_312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_167_ack_0, ack => inputPort_2_Daemon_CP_205_elements(47)); -- 
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/konst_169_sample_start__ps
      -- CP-element group 48: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/konst_169_sample_completed__ps
      -- CP-element group 48: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/konst_169_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/konst_169_sample_completed_
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/konst_169_update_start__ps
      -- CP-element group 49: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/konst_169_update_start_
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/konst_169_update_completed__ps
      -- 
    inputPort_2_Daemon_CP_205_elements(50) <= inputPort_2_Daemon_CP_205_elements(51);
    -- CP-element group 51:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	50 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/konst_169_update_completed_
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(51) is a control-delay.
    cp_element_51_delay: control_delay_element  generic map(name => " 51_delay", delay_value => 1)  port map(req => inputPort_2_Daemon_CP_205_elements(49), ack => inputPort_2_Daemon_CP_205_elements(51), clk => clk, reset =>reset);
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_Sample/req
      -- 
    req_333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(52), ack => next_last_dest_id_200_170_buf_req_0); -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_update_start_
      -- CP-element group 53: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_Update/req
      -- 
    req_338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(53), ack => next_last_dest_id_200_170_buf_req_1); -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_Sample/ack
      -- 
    ack_334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_200_170_buf_ack_0, ack => inputPort_2_Daemon_CP_205_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_Update/ack
      -- 
    ack_339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_200_170_buf_ack_1, ack => inputPort_2_Daemon_CP_205_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	42 
    -- CP-element group 56: 	38 
    -- CP-element group 56: 	20 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_1_212_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_1_212_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_1_212_Sample/req
      -- 
    req_348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(56), ack => WPIPE_noblock_obuf_2_1_212_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(42) & inputPort_2_Daemon_CP_205_elements(38) & inputPort_2_Daemon_CP_205_elements(20) & inputPort_2_Daemon_CP_205_elements(58);
      gj_inputPort_2_Daemon_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	40 
    -- CP-element group 57: 	34 
    -- CP-element group 57: 	16 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_1_212_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_1_212_update_start_
      -- CP-element group 57: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_1_212_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_1_212_Sample/ack
      -- CP-element group 57: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_1_212_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_1_212_Update/req
      -- 
    ack_349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_1_212_inst_ack_0, ack => inputPort_2_Daemon_CP_205_elements(57)); -- 
    req_353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(57), ack => WPIPE_noblock_obuf_2_1_212_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	69 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_1_212_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_1_212_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_1_212_Update/ack
      -- 
    ack_354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_1_212_inst_ack_1, ack => inputPort_2_Daemon_CP_205_elements(58)); -- 
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	42 
    -- CP-element group 59: 	38 
    -- CP-element group 59: 	20 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_2_221_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_2_221_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_2_221_Sample/req
      -- 
    req_362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(59), ack => WPIPE_noblock_obuf_2_2_221_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(42) & inputPort_2_Daemon_CP_205_elements(38) & inputPort_2_Daemon_CP_205_elements(20) & inputPort_2_Daemon_CP_205_elements(61);
      gj_inputPort_2_Daemon_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	40 
    -- CP-element group 60: 	34 
    -- CP-element group 60: 	16 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_2_221_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_2_221_update_start_
      -- CP-element group 60: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_2_221_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_2_221_Sample/ack
      -- CP-element group 60: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_2_221_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_2_221_Update/req
      -- 
    ack_363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_2_221_inst_ack_0, ack => inputPort_2_Daemon_CP_205_elements(60)); -- 
    req_367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(60), ack => WPIPE_noblock_obuf_2_2_221_inst_req_1); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	69 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_2_221_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_2_221_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_2_221_Update/ack
      -- 
    ack_368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_2_221_inst_ack_1, ack => inputPort_2_Daemon_CP_205_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	42 
    -- CP-element group 62: 	38 
    -- CP-element group 62: 	20 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_3_230_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_3_230_Sample/req
      -- CP-element group 62: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_3_230_sample_start_
      -- 
    req_376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(62), ack => WPIPE_noblock_obuf_2_3_230_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(42) & inputPort_2_Daemon_CP_205_elements(38) & inputPort_2_Daemon_CP_205_elements(20) & inputPort_2_Daemon_CP_205_elements(64);
      gj_inputPort_2_Daemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	40 
    -- CP-element group 63: 	34 
    -- CP-element group 63: 	16 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_3_230_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_3_230_Sample/ack
      -- CP-element group 63: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_3_230_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_3_230_Update/req
      -- CP-element group 63: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_3_230_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_3_230_update_start_
      -- 
    ack_377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_3_230_inst_ack_0, ack => inputPort_2_Daemon_CP_205_elements(63)); -- 
    req_381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(63), ack => WPIPE_noblock_obuf_2_3_230_inst_req_1); -- 
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	69 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_3_230_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_3_230_Update/ack
      -- CP-element group 64: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_3_230_update_completed_
      -- 
    ack_382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_3_230_inst_ack_1, ack => inputPort_2_Daemon_CP_205_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	42 
    -- CP-element group 65: 	38 
    -- CP-element group 65: 	20 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_4_239_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_4_239_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_4_239_Sample/req
      -- 
    req_390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(65), ack => WPIPE_noblock_obuf_2_4_239_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(42) & inputPort_2_Daemon_CP_205_elements(38) & inputPort_2_Daemon_CP_205_elements(20) & inputPort_2_Daemon_CP_205_elements(67);
      gj_inputPort_2_Daemon_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	40 
    -- CP-element group 66: 	34 
    -- CP-element group 66: 	16 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_4_239_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_4_239_update_start_
      -- CP-element group 66: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_4_239_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_4_239_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_4_239_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_4_239_Update/req
      -- 
    ack_391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_4_239_inst_ack_0, ack => inputPort_2_Daemon_CP_205_elements(66)); -- 
    req_395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(66), ack => WPIPE_noblock_obuf_2_4_239_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_4_239_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_4_239_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_4_239_Update/ack
      -- 
    ack_396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_4_239_inst_ack_1, ack => inputPort_2_Daemon_CP_205_elements(67)); -- 
    -- CP-element group 68:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	9 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	10 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(68) is a control-delay.
    cp_element_68_delay: control_delay_element  generic map(name => " 68_delay", delay_value => 1)  port map(req => inputPort_2_Daemon_CP_205_elements(9), ack => inputPort_2_Daemon_CP_205_elements(68), clk => clk, reset =>reset);
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	58 
    -- CP-element group 69: 	61 
    -- CP-element group 69: 	67 
    -- CP-element group 69: 	64 
    -- CP-element group 69: 	12 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	6 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/$exit
      -- 
    inputPort_2_Daemon_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(58) & inputPort_2_Daemon_CP_205_elements(61) & inputPort_2_Daemon_CP_205_elements(67) & inputPort_2_Daemon_CP_205_elements(64) & inputPort_2_Daemon_CP_205_elements(12);
      gj_inputPort_2_Daemon_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	5 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_156/do_while_stmt_157/loop_exit/$exit
      -- CP-element group 70: 	 branch_block_stmt_156/do_while_stmt_157/loop_exit/ack
      -- 
    ack_401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_157_branch_ack_0, ack => inputPort_2_Daemon_CP_205_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	5 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_156/do_while_stmt_157/loop_taken/$exit
      -- CP-element group 71: 	 branch_block_stmt_156/do_while_stmt_157/loop_taken/ack
      -- 
    ack_405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_157_branch_ack_1, ack => inputPort_2_Daemon_CP_205_elements(71)); -- 
    -- CP-element group 72:  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	3 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	1 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_156/do_while_stmt_157/$exit
      -- 
    inputPort_2_Daemon_CP_205_elements(72) <= inputPort_2_Daemon_CP_205_elements(3);
    inputPort_2_Daemon_do_while_stmt_157_terminator_406: loop_terminator -- 
      generic map (name => " inputPort_2_Daemon_do_while_stmt_157_terminator_406", max_iterations_in_flight =>7) 
      port map(loop_body_exit => inputPort_2_Daemon_CP_205_elements(6),loop_continue => inputPort_2_Daemon_CP_205_elements(71),loop_terminate => inputPort_2_Daemon_CP_205_elements(70),loop_back => inputPort_2_Daemon_CP_205_elements(4),loop_exit => inputPort_2_Daemon_CP_205_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_159_phi_seq_278_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_2_Daemon_CP_205_elements(21);
      inputPort_2_Daemon_CP_205_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_2_Daemon_CP_205_elements(28);
      inputPort_2_Daemon_CP_205_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_2_Daemon_CP_205_elements(29);
      inputPort_2_Daemon_CP_205_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_2_Daemon_CP_205_elements(23);
      inputPort_2_Daemon_CP_205_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_2_Daemon_CP_205_elements(30);
      inputPort_2_Daemon_CP_205_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_2_Daemon_CP_205_elements(32);
      inputPort_2_Daemon_CP_205_elements(24) <= phi_mux_reqs(1);
      phi_stmt_159_phi_seq_278 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_159_phi_seq_278") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_2_Daemon_CP_205_elements(17), 
          phi_sample_ack => inputPort_2_Daemon_CP_205_elements(18), 
          phi_update_req => inputPort_2_Daemon_CP_205_elements(19), 
          phi_update_ack => inputPort_2_Daemon_CP_205_elements(20), 
          phi_mux_ack => inputPort_2_Daemon_CP_205_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_167_phi_seq_340_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_2_Daemon_CP_205_elements(45);
      inputPort_2_Daemon_CP_205_elements(48)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_2_Daemon_CP_205_elements(48);
      inputPort_2_Daemon_CP_205_elements(49)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_2_Daemon_CP_205_elements(50);
      inputPort_2_Daemon_CP_205_elements(46) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_2_Daemon_CP_205_elements(43);
      inputPort_2_Daemon_CP_205_elements(52)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_2_Daemon_CP_205_elements(54);
      inputPort_2_Daemon_CP_205_elements(53)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_2_Daemon_CP_205_elements(55);
      inputPort_2_Daemon_CP_205_elements(44) <= phi_mux_reqs(1);
      phi_stmt_167_phi_seq_340 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_167_phi_seq_340") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_2_Daemon_CP_205_elements(11), 
          phi_sample_ack => inputPort_2_Daemon_CP_205_elements(41), 
          phi_update_req => inputPort_2_Daemon_CP_205_elements(13), 
          phi_update_ack => inputPort_2_Daemon_CP_205_elements(42), 
          phi_mux_ack => inputPort_2_Daemon_CP_205_elements(47), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_230_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= inputPort_2_Daemon_CP_205_elements(7);
        preds(1)  <= inputPort_2_Daemon_CP_205_elements(8);
        entry_tmerge_230 : transition_merge -- 
          generic map(name => " entry_tmerge_230")
          port map (preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal RPIPE_in_data_2_166_wire : std_logic_vector(31 downto 0);
    signal R_ONE_1_202_wire_constant : std_logic_vector(0 downto 0);
    signal SUB_u16_u16_189_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_192_wire : std_logic_vector(15 downto 0);
    signal count_down_159 : std_logic_vector(15 downto 0);
    signal data_to_outport_205 : std_logic_vector(32 downto 0);
    signal dest_id_180 : std_logic_vector(7 downto 0);
    signal input_word_164 : std_logic_vector(31 downto 0);
    signal konst_169_wire_constant : std_logic_vector(7 downto 0);
    signal konst_174_wire_constant : std_logic_vector(15 downto 0);
    signal konst_188_wire_constant : std_logic_vector(15 downto 0);
    signal konst_191_wire_constant : std_logic_vector(15 downto 0);
    signal konst_208_wire_constant : std_logic_vector(7 downto 0);
    signal konst_217_wire_constant : std_logic_vector(7 downto 0);
    signal konst_226_wire_constant : std_logic_vector(7 downto 0);
    signal konst_235_wire_constant : std_logic_vector(7 downto 0);
    signal konst_243_wire_constant : std_logic_vector(0 downto 0);
    signal last_dest_id_167 : std_logic_vector(7 downto 0);
    signal new_packet_176 : std_logic_vector(0 downto 0);
    signal next_count_down_194 : std_logic_vector(15 downto 0);
    signal next_count_down_194_161_buffered : std_logic_vector(15 downto 0);
    signal next_last_dest_id_200 : std_logic_vector(7 downto 0);
    signal next_last_dest_id_200_170_buffered : std_logic_vector(7 downto 0);
    signal pkt_length_184 : std_logic_vector(15 downto 0);
    signal send_to_1_210 : std_logic_vector(0 downto 0);
    signal send_to_2_219 : std_logic_vector(0 downto 0);
    signal send_to_3_228 : std_logic_vector(0 downto 0);
    signal send_to_4_237 : std_logic_vector(0 downto 0);
    signal type_cast_163_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    R_ONE_1_202_wire_constant <= "1";
    konst_169_wire_constant <= "00000000";
    konst_174_wire_constant <= "0000000000000000";
    konst_188_wire_constant <= "0000000000000001";
    konst_191_wire_constant <= "0000000000000001";
    konst_208_wire_constant <= "00000001";
    konst_217_wire_constant <= "00000010";
    konst_226_wire_constant <= "00000011";
    konst_235_wire_constant <= "00000100";
    konst_243_wire_constant <= "1";
    type_cast_163_wire_constant <= "0000000000000000";
    phi_stmt_159: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= next_count_down_194_161_buffered & type_cast_163_wire_constant;
      req <= phi_stmt_159_req_0 & phi_stmt_159_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_159",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_159_ack_0,
          idata => idata,
          odata => count_down_159,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_159
    phi_stmt_167: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_169_wire_constant & next_last_dest_id_200_170_buffered;
      req <= phi_stmt_167_req_0 & phi_stmt_167_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_167",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_167_ack_0,
          idata => idata,
          odata => last_dest_id_167,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_167
    -- flow-through select operator MUX_193_inst
    next_count_down_194 <= SUB_u16_u16_189_wire when (new_packet_176(0) /=  '0') else SUB_u16_u16_192_wire;
    -- flow-through select operator MUX_199_inst
    next_last_dest_id_200 <= dest_id_180 when (new_packet_176(0) /=  '0') else last_dest_id_167;
    -- flow-through slice operator slice_179_inst
    dest_id_180 <= input_word_164(31 downto 24);
    -- flow-through slice operator slice_183_inst
    pkt_length_184 <= input_word_164(23 downto 8);
    next_count_down_194_161_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_count_down_194_161_buf_req_0;
      next_count_down_194_161_buf_ack_0<= wack(0);
      rreq(0) <= next_count_down_194_161_buf_req_1;
      next_count_down_194_161_buf_ack_1<= rack(0);
      next_count_down_194_161_buf : InterlockBuffer generic map ( -- 
        name => "next_count_down_194_161_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_count_down_194,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_count_down_194_161_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_last_dest_id_200_170_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_last_dest_id_200_170_buf_req_0;
      next_last_dest_id_200_170_buf_ack_0<= wack(0);
      rreq(0) <= next_last_dest_id_200_170_buf_req_1;
      next_last_dest_id_200_170_buf_ack_1<= rack(0);
      next_last_dest_id_200_170_buf : InterlockBuffer generic map ( -- 
        name => "next_last_dest_id_200_170_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_last_dest_id_200,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_last_dest_id_200_170_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_164
    process(RPIPE_in_data_2_166_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := RPIPE_in_data_2_166_wire(31 downto 0);
      input_word_164 <= tmp_var; -- 
    end process;
    do_while_stmt_157_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_243_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_157_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_157_branch_req_0,
          ack0 => do_while_stmt_157_branch_ack_0,
          ack1 => do_while_stmt_157_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator CONCAT_u1_u33_204_inst
    process(R_ONE_1_202_wire_constant, input_word_164) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ONE_1_202_wire_constant, input_word_164, tmp_var);
      data_to_outport_205 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_175_inst
    process(count_down_159) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(count_down_159, konst_174_wire_constant, tmp_var);
      new_packet_176 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_209_inst
    process(next_last_dest_id_200) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_200, konst_208_wire_constant, tmp_var);
      send_to_1_210 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_218_inst
    process(next_last_dest_id_200) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_200, konst_217_wire_constant, tmp_var);
      send_to_2_219 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_227_inst
    process(next_last_dest_id_200) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_200, konst_226_wire_constant, tmp_var);
      send_to_3_228 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_236_inst
    process(next_last_dest_id_200) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_200, konst_235_wire_constant, tmp_var);
      send_to_4_237 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_189_inst
    process(pkt_length_184) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(pkt_length_184, konst_188_wire_constant, tmp_var);
      SUB_u16_u16_189_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_192_inst
    process(count_down_159) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(count_down_159, konst_191_wire_constant, tmp_var);
      SUB_u16_u16_192_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_in_data_2_166_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_in_data_2_166_inst_req_0;
      RPIPE_in_data_2_166_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_in_data_2_166_inst_req_1;
      RPIPE_in_data_2_166_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_in_data_2_166_wire <= data_out(31 downto 0);
      in_data_2_read_0_gI: SplitGuardInterface generic map(name => "in_data_2_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      in_data_2_read_0: InputPortRevised -- 
        generic map ( name => "in_data_2_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => in_data_2_pipe_read_req(0),
          oack => in_data_2_pipe_read_ack(0),
          odata => in_data_2_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_noblock_obuf_2_1_212_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_2_1_212_inst_req_0;
      WPIPE_noblock_obuf_2_1_212_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_2_1_212_inst_req_1;
      WPIPE_noblock_obuf_2_1_212_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_1_210(0);
      data_in <= data_to_outport_205;
      noblock_obuf_2_1_write_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_1_write_0: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_2_1", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_2_1_pipe_write_req(0),
          oack => noblock_obuf_2_1_pipe_write_ack(0),
          odata => noblock_obuf_2_1_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_noblock_obuf_2_2_221_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_2_2_221_inst_req_0;
      WPIPE_noblock_obuf_2_2_221_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_2_2_221_inst_req_1;
      WPIPE_noblock_obuf_2_2_221_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_2_219(0);
      data_in <= data_to_outport_205;
      noblock_obuf_2_2_write_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_2_write_1: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_2_2", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_2_2_pipe_write_req(0),
          oack => noblock_obuf_2_2_pipe_write_ack(0),
          odata => noblock_obuf_2_2_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_noblock_obuf_2_3_230_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_2_3_230_inst_req_0;
      WPIPE_noblock_obuf_2_3_230_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_2_3_230_inst_req_1;
      WPIPE_noblock_obuf_2_3_230_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_3_228(0);
      data_in <= data_to_outport_205;
      noblock_obuf_2_3_write_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_3_write_2: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_2_3", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_2_3_pipe_write_req(0),
          oack => noblock_obuf_2_3_pipe_write_ack(0),
          odata => noblock_obuf_2_3_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_noblock_obuf_2_4_239_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_2_4_239_inst_req_0;
      WPIPE_noblock_obuf_2_4_239_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_2_4_239_inst_req_1;
      WPIPE_noblock_obuf_2_4_239_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_4_237(0);
      data_in <= data_to_outport_205;
      noblock_obuf_2_4_write_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_4_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_4_write_3: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_2_4", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_2_4_pipe_write_req(0),
          oack => noblock_obuf_2_4_pipe_write_ack(0),
          odata => noblock_obuf_2_4_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end inputPort_2_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity inputPort_3_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    in_data_3_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_3_pipe_read_data : in   std_logic_vector(31 downto 0);
    noblock_obuf_3_2_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_2_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_3_3_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_3_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_3_4_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_4_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_3_1_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_1_pipe_write_data : out  std_logic_vector(32 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity inputPort_3_Daemon;
architecture inputPort_3_Daemon_arch of inputPort_3_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal inputPort_3_Daemon_CP_407_start: Boolean;
  signal inputPort_3_Daemon_CP_407_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_noblock_obuf_3_3_321_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_3_1_303_inst_ack_0 : boolean;
  signal next_count_down_285_254_buf_ack_1 : boolean;
  signal WPIPE_noblock_obuf_3_3_321_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_3_1_303_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_3_2_312_inst_req_1 : boolean;
  signal next_last_dest_id_291_261_buf_ack_1 : boolean;
  signal WPIPE_noblock_obuf_3_2_312_inst_ack_0 : boolean;
  signal next_count_down_285_254_buf_ack_0 : boolean;
  signal WPIPE_noblock_obuf_3_2_312_inst_req_0 : boolean;
  signal next_last_dest_id_291_261_buf_req_1 : boolean;
  signal next_count_down_285_254_buf_req_0 : boolean;
  signal next_count_down_285_254_buf_req_1 : boolean;
  signal WPIPE_noblock_obuf_3_4_330_inst_ack_1 : boolean;
  signal next_last_dest_id_291_261_buf_ack_0 : boolean;
  signal phi_stmt_258_req_0 : boolean;
  signal do_while_stmt_248_branch_req_0 : boolean;
  signal next_last_dest_id_291_261_buf_req_0 : boolean;
  signal WPIPE_noblock_obuf_3_3_321_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_3_4_330_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_3_3_321_inst_req_1 : boolean;
  signal do_while_stmt_248_branch_ack_1 : boolean;
  signal do_while_stmt_248_branch_ack_0 : boolean;
  signal phi_stmt_250_ack_0 : boolean;
  signal phi_stmt_250_req_0 : boolean;
  signal WPIPE_noblock_obuf_3_1_303_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_3_1_303_inst_req_1 : boolean;
  signal RPIPE_in_data_3_257_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_3_4_330_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_3_4_330_inst_req_0 : boolean;
  signal RPIPE_in_data_3_257_inst_req_1 : boolean;
  signal phi_stmt_258_req_1 : boolean;
  signal WPIPE_noblock_obuf_3_2_312_inst_ack_1 : boolean;
  signal RPIPE_in_data_3_257_inst_ack_0 : boolean;
  signal RPIPE_in_data_3_257_inst_req_0 : boolean;
  signal phi_stmt_258_ack_0 : boolean;
  signal phi_stmt_250_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "inputPort_3_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  inputPort_3_Daemon_CP_407_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "inputPort_3_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_3_Daemon_CP_407_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= inputPort_3_Daemon_CP_407_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_3_Daemon_CP_407_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  inputPort_3_Daemon_CP_407: Block -- control-path 
    signal inputPort_3_Daemon_CP_407_elements: BooleanArray(72 downto 0);
    -- 
  begin -- 
    inputPort_3_Daemon_CP_407_elements(0) <= inputPort_3_Daemon_CP_407_start;
    inputPort_3_Daemon_CP_407_symbol <= inputPort_3_Daemon_CP_407_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_247/$entry
      -- CP-element group 0: 	 branch_block_stmt_247/do_while_stmt_248__entry__
      -- CP-element group 0: 	 branch_block_stmt_247/branch_block_stmt_247__entry__
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	72 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_247/$exit
      -- CP-element group 1: 	 branch_block_stmt_247/do_while_stmt_248__exit__
      -- CP-element group 1: 	 branch_block_stmt_247/branch_block_stmt_247__exit__
      -- CP-element group 1: 	 $exit
      -- 
    inputPort_3_Daemon_CP_407_elements(1) <= inputPort_3_Daemon_CP_407_elements(72);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248__entry__
      -- CP-element group 2: 	 branch_block_stmt_247/do_while_stmt_248/$entry
      -- 
    inputPort_3_Daemon_CP_407_elements(2) <= inputPort_3_Daemon_CP_407_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	72 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248__exit__
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_247/do_while_stmt_248/loop_back
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	71 
    -- CP-element group 5: 	70 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_247/do_while_stmt_248/condition_done
      -- CP-element group 5: 	 branch_block_stmt_247/do_while_stmt_248/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_247/do_while_stmt_248/loop_exit/$entry
      -- 
    inputPort_3_Daemon_CP_407_elements(5) <= inputPort_3_Daemon_CP_407_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	69 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_247/do_while_stmt_248/loop_body_done
      -- 
    inputPort_3_Daemon_CP_407_elements(6) <= inputPort_3_Daemon_CP_407_elements(69);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	43 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/back_edge_to_loop_body
      -- 
    inputPort_3_Daemon_CP_407_elements(7) <= inputPort_3_Daemon_CP_407_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	45 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/first_time_through_loop_body
      -- 
    inputPort_3_Daemon_CP_407_elements(8) <= inputPort_3_Daemon_CP_407_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	37 
    -- CP-element group 9: 	38 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	68 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_255_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/$entry
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	68 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/condition_evaluated
      -- 
    condition_evaluated_431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(10), ack => do_while_stmt_248_branch_req_0); -- 
    inputPort_3_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(14) & inputPort_3_Daemon_CP_407_elements(68);
      gj_inputPort_3_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	37 
    -- CP-element group 11: 	9 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	39 
    -- CP-element group 11: 	33 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_sample_start__ps
      -- 
    inputPort_3_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(15) & inputPort_3_Daemon_CP_407_elements(37) & inputPort_3_Daemon_CP_407_elements(9) & inputPort_3_Daemon_CP_407_elements(14);
      gj_inputPort_3_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	40 
    -- CP-element group 12: 	35 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	69 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	37 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_255_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_sample_completed_
      -- 
    inputPort_3_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(17) & inputPort_3_Daemon_CP_407_elements(40) & inputPort_3_Daemon_CP_407_elements(35);
      gj_inputPort_3_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	38 
    -- CP-element group 13: 	32 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	41 
    -- CP-element group 13: 	34 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_update_start__ps
      -- 
    inputPort_3_Daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(16) & inputPort_3_Daemon_CP_407_elements(38) & inputPort_3_Daemon_CP_407_elements(32);
      gj_inputPort_3_Daemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	42 
    -- CP-element group 14: 	36 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/aggregated_phi_update_ack
      -- 
    inputPort_3_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(18) & inputPort_3_Daemon_CP_407_elements(42) & inputPort_3_Daemon_CP_407_elements(36);
      gj_inputPort_3_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_sample_start_
      -- 
    inputPort_3_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(9) & inputPort_3_Daemon_CP_407_elements(12);
      gj_inputPort_3_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	57 
    -- CP-element group 16: 	60 
    -- CP-element group 16: 	63 
    -- CP-element group 16: 	66 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_update_start_
      -- 
    inputPort_3_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(9) & inputPort_3_Daemon_CP_407_elements(57) & inputPort_3_Daemon_CP_407_elements(60) & inputPort_3_Daemon_CP_407_elements(63) & inputPort_3_Daemon_CP_407_elements(66);
      gj_inputPort_3_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_sample_completed__ps
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	56 
    -- CP-element group 18: 	59 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	62 
    -- CP-element group 18: 	65 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_update_completed_
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_loopback_trigger
      -- 
    inputPort_3_Daemon_CP_407_elements(19) <= inputPort_3_Daemon_CP_407_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_loopback_sample_req_ps
      -- CP-element group 20: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_loopback_sample_req
      -- 
    phi_stmt_250_loopback_sample_req_446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_250_loopback_sample_req_446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(20), ack => phi_stmt_250_req_1); -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_entry_trigger
      -- 
    inputPort_3_Daemon_CP_407_elements(21) <= inputPort_3_Daemon_CP_407_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_entry_sample_req_ps
      -- CP-element group 22: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_entry_sample_req
      -- 
    phi_stmt_250_entry_sample_req_449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_250_entry_sample_req_449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(22), ack => phi_stmt_250_req_0); -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_phi_mux_ack_ps
      -- CP-element group 23: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_phi_mux_ack
      -- 
    phi_stmt_250_phi_mux_ack_452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_250_ack_0, ack => inputPort_3_Daemon_CP_407_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/type_cast_253_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/type_cast_253_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/type_cast_253_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/type_cast_253_sample_start__ps
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/type_cast_253_update_start_
      -- CP-element group 25: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/type_cast_253_update_start__ps
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/type_cast_253_update_completed__ps
      -- 
    inputPort_3_Daemon_CP_407_elements(26) <= inputPort_3_Daemon_CP_407_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/type_cast_253_update_completed_
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => inputPort_3_Daemon_CP_407_elements(25), ack => inputPort_3_Daemon_CP_407_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_Sample/req
      -- CP-element group 28: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_sample_start__ps
      -- 
    req_473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(28), ack => next_count_down_285_254_buf_req_0); -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_Update/req
      -- CP-element group 29: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_update_start_
      -- CP-element group 29: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_update_start__ps
      -- 
    req_478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(29), ack => next_count_down_285_254_buf_req_1); -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_Sample/ack
      -- CP-element group 30: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_sample_completed__ps
      -- 
    ack_474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_285_254_buf_ack_0, ack => inputPort_3_Daemon_CP_407_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_Update/ack
      -- CP-element group 31: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_update_completed__ps
      -- 
    ack_479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_285_254_buf_ack_1, ack => inputPort_3_Daemon_CP_407_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	57 
    -- CP-element group 32: 	60 
    -- CP-element group 32: 	63 
    -- CP-element group 32: 	66 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_255_update_start_
      -- 
    inputPort_3_Daemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(9) & inputPort_3_Daemon_CP_407_elements(57) & inputPort_3_Daemon_CP_407_elements(60) & inputPort_3_Daemon_CP_407_elements(63) & inputPort_3_Daemon_CP_407_elements(66);
      gj_inputPort_3_Daemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/RPIPE_in_data_3_257_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/RPIPE_in_data_3_257_Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/RPIPE_in_data_3_257_Sample/$entry
      -- 
    rr_492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(33), ack => RPIPE_in_data_3_257_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(11) & inputPort_3_Daemon_CP_407_elements(36);
      gj_inputPort_3_Daemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	13 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/RPIPE_in_data_3_257_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/RPIPE_in_data_3_257_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/RPIPE_in_data_3_257_update_start_
      -- 
    cr_497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(34), ack => RPIPE_in_data_3_257_inst_req_1); -- 
    inputPort_3_Daemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(35) & inputPort_3_Daemon_CP_407_elements(13);
      gj_inputPort_3_Daemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: 	12 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/RPIPE_in_data_3_257_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/RPIPE_in_data_3_257_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/RPIPE_in_data_3_257_Sample/$exit
      -- 
    ra_493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_3_257_inst_ack_0, ack => inputPort_3_Daemon_CP_407_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	56 
    -- CP-element group 36: 	59 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	62 
    -- CP-element group 36: 	65 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_255_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/RPIPE_in_data_3_257_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/RPIPE_in_data_3_257_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/RPIPE_in_data_3_257_update_completed_
      -- 
    ca_498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_3_257_inst_ack_1, ack => inputPort_3_Daemon_CP_407_elements(36)); -- 
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	9 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	12 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	11 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_sample_start_
      -- 
    inputPort_3_Daemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(9) & inputPort_3_Daemon_CP_407_elements(12);
      gj_inputPort_3_Daemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	9 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	57 
    -- CP-element group 38: 	60 
    -- CP-element group 38: 	63 
    -- CP-element group 38: 	66 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	13 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_update_start_
      -- 
    inputPort_3_Daemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(9) & inputPort_3_Daemon_CP_407_elements(57) & inputPort_3_Daemon_CP_407_elements(60) & inputPort_3_Daemon_CP_407_elements(63) & inputPort_3_Daemon_CP_407_elements(66);
      gj_inputPort_3_Daemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	11 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_sample_start__ps
      -- 
    inputPort_3_Daemon_CP_407_elements(39) <= inputPort_3_Daemon_CP_407_elements(11);
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	12 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_sample_completed__ps
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	13 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_update_start__ps
      -- 
    inputPort_3_Daemon_CP_407_elements(41) <= inputPort_3_Daemon_CP_407_elements(13);
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	56 
    -- CP-element group 42: 	59 
    -- CP-element group 42: 	14 
    -- CP-element group 42: 	62 
    -- CP-element group 42: 	65 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_update_completed__ps
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	7 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_loopback_trigger
      -- 
    inputPort_3_Daemon_CP_407_elements(43) <= inputPort_3_Daemon_CP_407_elements(7);
    -- CP-element group 44:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_loopback_sample_req_ps
      -- CP-element group 44: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_loopback_sample_req
      -- 
    phi_stmt_258_loopback_sample_req_508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_258_loopback_sample_req_508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(44), ack => phi_stmt_258_req_1); -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	8 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_entry_trigger
      -- 
    inputPort_3_Daemon_CP_407_elements(45) <= inputPort_3_Daemon_CP_407_elements(8);
    -- CP-element group 46:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_entry_sample_req_ps
      -- CP-element group 46: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_entry_sample_req
      -- 
    phi_stmt_258_entry_sample_req_511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_258_entry_sample_req_511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(46), ack => phi_stmt_258_req_0); -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_phi_mux_ack_ps
      -- CP-element group 47: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_phi_mux_ack
      -- 
    phi_stmt_258_phi_mux_ack_514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_258_ack_0, ack => inputPort_3_Daemon_CP_407_elements(47)); -- 
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/konst_260_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/konst_260_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/konst_260_sample_completed__ps
      -- CP-element group 48: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/konst_260_sample_start__ps
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/konst_260_update_start__ps
      -- CP-element group 49: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/konst_260_update_start_
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/konst_260_update_completed__ps
      -- 
    inputPort_3_Daemon_CP_407_elements(50) <= inputPort_3_Daemon_CP_407_elements(51);
    -- CP-element group 51:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	50 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/konst_260_update_completed_
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(51) is a control-delay.
    cp_element_51_delay: control_delay_element  generic map(name => " 51_delay", delay_value => 1)  port map(req => inputPort_3_Daemon_CP_407_elements(49), ack => inputPort_3_Daemon_CP_407_elements(51), clk => clk, reset =>reset);
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_Sample/req
      -- CP-element group 52: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_sample_start__ps
      -- 
    req_535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(52), ack => next_last_dest_id_291_261_buf_req_0); -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_Update/req
      -- CP-element group 53: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_update_start_
      -- CP-element group 53: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_update_start__ps
      -- 
    req_540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(53), ack => next_last_dest_id_291_261_buf_req_1); -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_Sample/ack
      -- CP-element group 54: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_sample_completed__ps
      -- 
    ack_536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_291_261_buf_ack_0, ack => inputPort_3_Daemon_CP_407_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_Update/ack
      -- CP-element group 55: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_update_completed__ps
      -- 
    ack_541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_291_261_buf_ack_1, ack => inputPort_3_Daemon_CP_407_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	18 
    -- CP-element group 56: 	42 
    -- CP-element group 56: 	36 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_1_303_Sample/req
      -- CP-element group 56: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_1_303_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_1_303_sample_start_
      -- 
    req_550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(56), ack => WPIPE_noblock_obuf_3_1_303_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 7,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(18) & inputPort_3_Daemon_CP_407_elements(42) & inputPort_3_Daemon_CP_407_elements(36) & inputPort_3_Daemon_CP_407_elements(58);
      gj_inputPort_3_Daemon_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	16 
    -- CP-element group 57: 	38 
    -- CP-element group 57: 	32 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_1_303_Sample/ack
      -- CP-element group 57: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_1_303_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_1_303_update_start_
      -- CP-element group 57: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_1_303_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_1_303_Update/req
      -- CP-element group 57: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_1_303_Update/$entry
      -- 
    ack_551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_1_303_inst_ack_0, ack => inputPort_3_Daemon_CP_407_elements(57)); -- 
    req_555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(57), ack => WPIPE_noblock_obuf_3_1_303_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	69 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_1_303_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_1_303_Update/ack
      -- CP-element group 58: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_1_303_Update/$exit
      -- 
    ack_556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_1_303_inst_ack_1, ack => inputPort_3_Daemon_CP_407_elements(58)); -- 
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	18 
    -- CP-element group 59: 	42 
    -- CP-element group 59: 	36 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_2_312_Sample/req
      -- CP-element group 59: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_2_312_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_2_312_sample_start_
      -- 
    req_564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(59), ack => WPIPE_noblock_obuf_3_2_312_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 7,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(18) & inputPort_3_Daemon_CP_407_elements(42) & inputPort_3_Daemon_CP_407_elements(36) & inputPort_3_Daemon_CP_407_elements(61);
      gj_inputPort_3_Daemon_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	16 
    -- CP-element group 60: 	38 
    -- CP-element group 60: 	32 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_2_312_Update/req
      -- CP-element group 60: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_2_312_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_2_312_Sample/ack
      -- CP-element group 60: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_2_312_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_2_312_update_start_
      -- CP-element group 60: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_2_312_sample_completed_
      -- 
    ack_565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_2_312_inst_ack_0, ack => inputPort_3_Daemon_CP_407_elements(60)); -- 
    req_569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(60), ack => WPIPE_noblock_obuf_3_2_312_inst_req_1); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	69 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_2_312_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_2_312_Update/ack
      -- CP-element group 61: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_2_312_update_completed_
      -- 
    ack_570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_2_312_inst_ack_1, ack => inputPort_3_Daemon_CP_407_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	18 
    -- CP-element group 62: 	42 
    -- CP-element group 62: 	36 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_3_321_Sample/req
      -- CP-element group 62: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_3_321_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_3_321_sample_start_
      -- 
    req_578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(62), ack => WPIPE_noblock_obuf_3_3_321_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 7,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(18) & inputPort_3_Daemon_CP_407_elements(42) & inputPort_3_Daemon_CP_407_elements(36) & inputPort_3_Daemon_CP_407_elements(64);
      gj_inputPort_3_Daemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	16 
    -- CP-element group 63: 	38 
    -- CP-element group 63: 	32 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_3_321_Sample/ack
      -- CP-element group 63: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_3_321_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_3_321_Update/req
      -- CP-element group 63: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_3_321_update_start_
      -- CP-element group 63: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_3_321_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_3_321_Update/$entry
      -- 
    ack_579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_3_321_inst_ack_0, ack => inputPort_3_Daemon_CP_407_elements(63)); -- 
    req_583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(63), ack => WPIPE_noblock_obuf_3_3_321_inst_req_1); -- 
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	69 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_3_321_Update/ack
      -- CP-element group 64: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_3_321_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_3_321_Update/$exit
      -- 
    ack_584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_3_321_inst_ack_1, ack => inputPort_3_Daemon_CP_407_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	18 
    -- CP-element group 65: 	42 
    -- CP-element group 65: 	36 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_4_330_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_4_330_Sample/req
      -- CP-element group 65: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_4_330_Sample/$entry
      -- 
    req_592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(65), ack => WPIPE_noblock_obuf_3_4_330_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 7,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(18) & inputPort_3_Daemon_CP_407_elements(42) & inputPort_3_Daemon_CP_407_elements(36) & inputPort_3_Daemon_CP_407_elements(67);
      gj_inputPort_3_Daemon_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	16 
    -- CP-element group 66: 	38 
    -- CP-element group 66: 	32 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_4_330_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_4_330_Update/req
      -- CP-element group 66: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_4_330_update_start_
      -- CP-element group 66: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_4_330_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_4_330_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_4_330_Sample/$exit
      -- 
    ack_593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_4_330_inst_ack_0, ack => inputPort_3_Daemon_CP_407_elements(66)); -- 
    req_597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(66), ack => WPIPE_noblock_obuf_3_4_330_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_4_330_Update/ack
      -- CP-element group 67: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_4_330_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_4_330_update_completed_
      -- 
    ack_598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_4_330_inst_ack_1, ack => inputPort_3_Daemon_CP_407_elements(67)); -- 
    -- CP-element group 68:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	9 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	10 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(68) is a control-delay.
    cp_element_68_delay: control_delay_element  generic map(name => " 68_delay", delay_value => 1)  port map(req => inputPort_3_Daemon_CP_407_elements(9), ack => inputPort_3_Daemon_CP_407_elements(68), clk => clk, reset =>reset);
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	58 
    -- CP-element group 69: 	12 
    -- CP-element group 69: 	61 
    -- CP-element group 69: 	64 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	6 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/$exit
      -- 
    inputPort_3_Daemon_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(58) & inputPort_3_Daemon_CP_407_elements(12) & inputPort_3_Daemon_CP_407_elements(61) & inputPort_3_Daemon_CP_407_elements(64) & inputPort_3_Daemon_CP_407_elements(67);
      gj_inputPort_3_Daemon_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	5 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_247/do_while_stmt_248/loop_exit/ack
      -- CP-element group 70: 	 branch_block_stmt_247/do_while_stmt_248/loop_exit/$exit
      -- 
    ack_603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_248_branch_ack_0, ack => inputPort_3_Daemon_CP_407_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	5 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_247/do_while_stmt_248/loop_taken/ack
      -- CP-element group 71: 	 branch_block_stmt_247/do_while_stmt_248/loop_taken/$exit
      -- 
    ack_607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_248_branch_ack_1, ack => inputPort_3_Daemon_CP_407_elements(71)); -- 
    -- CP-element group 72:  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	3 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	1 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_247/do_while_stmt_248/$exit
      -- 
    inputPort_3_Daemon_CP_407_elements(72) <= inputPort_3_Daemon_CP_407_elements(3);
    inputPort_3_Daemon_do_while_stmt_248_terminator_608: loop_terminator -- 
      generic map (name => " inputPort_3_Daemon_do_while_stmt_248_terminator_608", max_iterations_in_flight =>7) 
      port map(loop_body_exit => inputPort_3_Daemon_CP_407_elements(6),loop_continue => inputPort_3_Daemon_CP_407_elements(71),loop_terminate => inputPort_3_Daemon_CP_407_elements(70),loop_back => inputPort_3_Daemon_CP_407_elements(4),loop_exit => inputPort_3_Daemon_CP_407_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_250_phi_seq_480_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_3_Daemon_CP_407_elements(21);
      inputPort_3_Daemon_CP_407_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_3_Daemon_CP_407_elements(24);
      inputPort_3_Daemon_CP_407_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_3_Daemon_CP_407_elements(26);
      inputPort_3_Daemon_CP_407_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_3_Daemon_CP_407_elements(19);
      inputPort_3_Daemon_CP_407_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_3_Daemon_CP_407_elements(30);
      inputPort_3_Daemon_CP_407_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_3_Daemon_CP_407_elements(31);
      inputPort_3_Daemon_CP_407_elements(20) <= phi_mux_reqs(1);
      phi_stmt_250_phi_seq_480 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_250_phi_seq_480") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_3_Daemon_CP_407_elements(11), 
          phi_sample_ack => inputPort_3_Daemon_CP_407_elements(17), 
          phi_update_req => inputPort_3_Daemon_CP_407_elements(13), 
          phi_update_ack => inputPort_3_Daemon_CP_407_elements(18), 
          phi_mux_ack => inputPort_3_Daemon_CP_407_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_258_phi_seq_542_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_3_Daemon_CP_407_elements(45);
      inputPort_3_Daemon_CP_407_elements(48)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_3_Daemon_CP_407_elements(48);
      inputPort_3_Daemon_CP_407_elements(49)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_3_Daemon_CP_407_elements(50);
      inputPort_3_Daemon_CP_407_elements(46) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_3_Daemon_CP_407_elements(43);
      inputPort_3_Daemon_CP_407_elements(52)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_3_Daemon_CP_407_elements(54);
      inputPort_3_Daemon_CP_407_elements(53)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_3_Daemon_CP_407_elements(55);
      inputPort_3_Daemon_CP_407_elements(44) <= phi_mux_reqs(1);
      phi_stmt_258_phi_seq_542 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_258_phi_seq_542") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_3_Daemon_CP_407_elements(39), 
          phi_sample_ack => inputPort_3_Daemon_CP_407_elements(40), 
          phi_update_req => inputPort_3_Daemon_CP_407_elements(41), 
          phi_update_ack => inputPort_3_Daemon_CP_407_elements(42), 
          phi_mux_ack => inputPort_3_Daemon_CP_407_elements(47), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_432_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= inputPort_3_Daemon_CP_407_elements(7);
        preds(1)  <= inputPort_3_Daemon_CP_407_elements(8);
        entry_tmerge_432 : transition_merge -- 
          generic map(name => " entry_tmerge_432")
          port map (preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal RPIPE_in_data_3_257_wire : std_logic_vector(31 downto 0);
    signal R_ONE_1_293_wire_constant : std_logic_vector(0 downto 0);
    signal SUB_u16_u16_280_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_283_wire : std_logic_vector(15 downto 0);
    signal count_down_250 : std_logic_vector(15 downto 0);
    signal data_to_outport_296 : std_logic_vector(32 downto 0);
    signal dest_id_271 : std_logic_vector(7 downto 0);
    signal input_word_255 : std_logic_vector(31 downto 0);
    signal konst_260_wire_constant : std_logic_vector(7 downto 0);
    signal konst_265_wire_constant : std_logic_vector(15 downto 0);
    signal konst_279_wire_constant : std_logic_vector(15 downto 0);
    signal konst_282_wire_constant : std_logic_vector(15 downto 0);
    signal konst_299_wire_constant : std_logic_vector(7 downto 0);
    signal konst_308_wire_constant : std_logic_vector(7 downto 0);
    signal konst_317_wire_constant : std_logic_vector(7 downto 0);
    signal konst_326_wire_constant : std_logic_vector(7 downto 0);
    signal konst_334_wire_constant : std_logic_vector(0 downto 0);
    signal last_dest_id_258 : std_logic_vector(7 downto 0);
    signal new_packet_267 : std_logic_vector(0 downto 0);
    signal next_count_down_285 : std_logic_vector(15 downto 0);
    signal next_count_down_285_254_buffered : std_logic_vector(15 downto 0);
    signal next_last_dest_id_291 : std_logic_vector(7 downto 0);
    signal next_last_dest_id_291_261_buffered : std_logic_vector(7 downto 0);
    signal pkt_length_275 : std_logic_vector(15 downto 0);
    signal send_to_1_301 : std_logic_vector(0 downto 0);
    signal send_to_2_310 : std_logic_vector(0 downto 0);
    signal send_to_3_319 : std_logic_vector(0 downto 0);
    signal send_to_4_328 : std_logic_vector(0 downto 0);
    signal type_cast_253_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    R_ONE_1_293_wire_constant <= "1";
    konst_260_wire_constant <= "00000000";
    konst_265_wire_constant <= "0000000000000000";
    konst_279_wire_constant <= "0000000000000001";
    konst_282_wire_constant <= "0000000000000001";
    konst_299_wire_constant <= "00000001";
    konst_308_wire_constant <= "00000010";
    konst_317_wire_constant <= "00000011";
    konst_326_wire_constant <= "00000100";
    konst_334_wire_constant <= "1";
    type_cast_253_wire_constant <= "0000000000000000";
    phi_stmt_250: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_253_wire_constant & next_count_down_285_254_buffered;
      req <= phi_stmt_250_req_0 & phi_stmt_250_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_250",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_250_ack_0,
          idata => idata,
          odata => count_down_250,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_250
    phi_stmt_258: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_260_wire_constant & next_last_dest_id_291_261_buffered;
      req <= phi_stmt_258_req_0 & phi_stmt_258_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_258",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_258_ack_0,
          idata => idata,
          odata => last_dest_id_258,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_258
    -- flow-through select operator MUX_284_inst
    next_count_down_285 <= SUB_u16_u16_280_wire when (new_packet_267(0) /=  '0') else SUB_u16_u16_283_wire;
    -- flow-through select operator MUX_290_inst
    next_last_dest_id_291 <= dest_id_271 when (new_packet_267(0) /=  '0') else last_dest_id_258;
    -- flow-through slice operator slice_270_inst
    dest_id_271 <= input_word_255(31 downto 24);
    -- flow-through slice operator slice_274_inst
    pkt_length_275 <= input_word_255(23 downto 8);
    next_count_down_285_254_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_count_down_285_254_buf_req_0;
      next_count_down_285_254_buf_ack_0<= wack(0);
      rreq(0) <= next_count_down_285_254_buf_req_1;
      next_count_down_285_254_buf_ack_1<= rack(0);
      next_count_down_285_254_buf : InterlockBuffer generic map ( -- 
        name => "next_count_down_285_254_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_count_down_285,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_count_down_285_254_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_last_dest_id_291_261_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_last_dest_id_291_261_buf_req_0;
      next_last_dest_id_291_261_buf_ack_0<= wack(0);
      rreq(0) <= next_last_dest_id_291_261_buf_req_1;
      next_last_dest_id_291_261_buf_ack_1<= rack(0);
      next_last_dest_id_291_261_buf : InterlockBuffer generic map ( -- 
        name => "next_last_dest_id_291_261_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_last_dest_id_291,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_last_dest_id_291_261_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_255
    process(RPIPE_in_data_3_257_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := RPIPE_in_data_3_257_wire(31 downto 0);
      input_word_255 <= tmp_var; -- 
    end process;
    do_while_stmt_248_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_334_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_248_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_248_branch_req_0,
          ack0 => do_while_stmt_248_branch_ack_0,
          ack1 => do_while_stmt_248_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator CONCAT_u1_u33_295_inst
    process(R_ONE_1_293_wire_constant, input_word_255) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ONE_1_293_wire_constant, input_word_255, tmp_var);
      data_to_outport_296 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_266_inst
    process(count_down_250) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(count_down_250, konst_265_wire_constant, tmp_var);
      new_packet_267 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_300_inst
    process(next_last_dest_id_291) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_291, konst_299_wire_constant, tmp_var);
      send_to_1_301 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_309_inst
    process(next_last_dest_id_291) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_291, konst_308_wire_constant, tmp_var);
      send_to_2_310 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_318_inst
    process(next_last_dest_id_291) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_291, konst_317_wire_constant, tmp_var);
      send_to_3_319 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_327_inst
    process(next_last_dest_id_291) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_291, konst_326_wire_constant, tmp_var);
      send_to_4_328 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_280_inst
    process(pkt_length_275) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(pkt_length_275, konst_279_wire_constant, tmp_var);
      SUB_u16_u16_280_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_283_inst
    process(count_down_250) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(count_down_250, konst_282_wire_constant, tmp_var);
      SUB_u16_u16_283_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_in_data_3_257_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_in_data_3_257_inst_req_0;
      RPIPE_in_data_3_257_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_in_data_3_257_inst_req_1;
      RPIPE_in_data_3_257_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_in_data_3_257_wire <= data_out(31 downto 0);
      in_data_3_read_0_gI: SplitGuardInterface generic map(name => "in_data_3_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      in_data_3_read_0: InputPortRevised -- 
        generic map ( name => "in_data_3_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => in_data_3_pipe_read_req(0),
          oack => in_data_3_pipe_read_ack(0),
          odata => in_data_3_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_noblock_obuf_3_1_303_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_3_1_303_inst_req_0;
      WPIPE_noblock_obuf_3_1_303_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_3_1_303_inst_req_1;
      WPIPE_noblock_obuf_3_1_303_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_1_301(0);
      data_in <= data_to_outport_296;
      noblock_obuf_3_1_write_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_1_write_0: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_3_1", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_3_1_pipe_write_req(0),
          oack => noblock_obuf_3_1_pipe_write_ack(0),
          odata => noblock_obuf_3_1_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_noblock_obuf_3_2_312_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_3_2_312_inst_req_0;
      WPIPE_noblock_obuf_3_2_312_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_3_2_312_inst_req_1;
      WPIPE_noblock_obuf_3_2_312_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_2_310(0);
      data_in <= data_to_outport_296;
      noblock_obuf_3_2_write_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_2_write_1: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_3_2", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_3_2_pipe_write_req(0),
          oack => noblock_obuf_3_2_pipe_write_ack(0),
          odata => noblock_obuf_3_2_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_noblock_obuf_3_3_321_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_3_3_321_inst_req_0;
      WPIPE_noblock_obuf_3_3_321_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_3_3_321_inst_req_1;
      WPIPE_noblock_obuf_3_3_321_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_3_319(0);
      data_in <= data_to_outport_296;
      noblock_obuf_3_3_write_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_3_write_2: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_3_3", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_3_3_pipe_write_req(0),
          oack => noblock_obuf_3_3_pipe_write_ack(0),
          odata => noblock_obuf_3_3_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_noblock_obuf_3_4_330_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_3_4_330_inst_req_0;
      WPIPE_noblock_obuf_3_4_330_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_3_4_330_inst_req_1;
      WPIPE_noblock_obuf_3_4_330_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_4_328(0);
      data_in <= data_to_outport_296;
      noblock_obuf_3_4_write_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_4_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_4_write_3: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_3_4", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_3_4_pipe_write_req(0),
          oack => noblock_obuf_3_4_pipe_write_ack(0),
          odata => noblock_obuf_3_4_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end inputPort_3_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity inputPort_4_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    in_data_4_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_4_pipe_read_data : in   std_logic_vector(31 downto 0);
    noblock_obuf_4_1_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_1_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_4_2_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_2_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_4_3_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_3_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_4_4_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_4_pipe_write_data : out  std_logic_vector(32 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity inputPort_4_Daemon;
architecture inputPort_4_Daemon_arch of inputPort_4_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal inputPort_4_Daemon_CP_609_start: Boolean;
  signal inputPort_4_Daemon_CP_609_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_339_branch_req_0 : boolean;
  signal phi_stmt_341_req_1 : boolean;
  signal phi_stmt_341_req_0 : boolean;
  signal phi_stmt_341_ack_0 : boolean;
  signal next_count_down_376_345_buf_req_0 : boolean;
  signal next_count_down_376_345_buf_ack_0 : boolean;
  signal next_count_down_376_345_buf_req_1 : boolean;
  signal next_count_down_376_345_buf_ack_1 : boolean;
  signal RPIPE_in_data_4_348_inst_req_0 : boolean;
  signal RPIPE_in_data_4_348_inst_ack_0 : boolean;
  signal RPIPE_in_data_4_348_inst_req_1 : boolean;
  signal RPIPE_in_data_4_348_inst_ack_1 : boolean;
  signal phi_stmt_349_req_1 : boolean;
  signal phi_stmt_349_req_0 : boolean;
  signal phi_stmt_349_ack_0 : boolean;
  signal next_last_dest_id_382_352_buf_req_0 : boolean;
  signal next_last_dest_id_382_352_buf_ack_0 : boolean;
  signal next_last_dest_id_382_352_buf_req_1 : boolean;
  signal next_last_dest_id_382_352_buf_ack_1 : boolean;
  signal WPIPE_noblock_obuf_4_1_394_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_4_1_394_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_4_1_394_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_4_1_394_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_4_2_403_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_4_2_403_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_4_2_403_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_4_2_403_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_4_3_412_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_4_3_412_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_4_3_412_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_4_3_412_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_4_4_421_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_4_4_421_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_4_4_421_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_4_4_421_inst_ack_1 : boolean;
  signal do_while_stmt_339_branch_ack_0 : boolean;
  signal do_while_stmt_339_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "inputPort_4_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  inputPort_4_Daemon_CP_609_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "inputPort_4_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_4_Daemon_CP_609_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= inputPort_4_Daemon_CP_609_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_4_Daemon_CP_609_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  inputPort_4_Daemon_CP_609: Block -- control-path 
    signal inputPort_4_Daemon_CP_609_elements: BooleanArray(72 downto 0);
    -- 
  begin -- 
    inputPort_4_Daemon_CP_609_elements(0) <= inputPort_4_Daemon_CP_609_start;
    inputPort_4_Daemon_CP_609_symbol <= inputPort_4_Daemon_CP_609_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_338/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_338/branch_block_stmt_338__entry__
      -- CP-element group 0: 	 branch_block_stmt_338/do_while_stmt_339__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	72 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_338/branch_block_stmt_338__exit__
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_338/$exit
      -- CP-element group 1: 	 branch_block_stmt_338/do_while_stmt_339__exit__
      -- 
    inputPort_4_Daemon_CP_609_elements(1) <= inputPort_4_Daemon_CP_609_elements(72);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_338/do_while_stmt_339/$entry
      -- CP-element group 2: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339__entry__
      -- 
    inputPort_4_Daemon_CP_609_elements(2) <= inputPort_4_Daemon_CP_609_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	72 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339__exit__
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_338/do_while_stmt_339/loop_back
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	70 
    -- CP-element group 5: 	71 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_338/do_while_stmt_339/condition_done
      -- CP-element group 5: 	 branch_block_stmt_338/do_while_stmt_339/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_338/do_while_stmt_339/loop_taken/$entry
      -- 
    inputPort_4_Daemon_CP_609_elements(5) <= inputPort_4_Daemon_CP_609_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	69 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_338/do_while_stmt_339/loop_body_done
      -- 
    inputPort_4_Daemon_CP_609_elements(6) <= inputPort_4_Daemon_CP_609_elements(69);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	43 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/back_edge_to_loop_body
      -- 
    inputPort_4_Daemon_CP_609_elements(7) <= inputPort_4_Daemon_CP_609_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	45 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/first_time_through_loop_body
      -- 
    inputPort_4_Daemon_CP_609_elements(8) <= inputPort_4_Daemon_CP_609_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	37 
    -- CP-element group 9: 	38 
    -- CP-element group 9: 	68 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_346_sample_start_
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	68 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/condition_evaluated
      -- 
    condition_evaluated_633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(10), ack => do_while_stmt_339_branch_req_0); -- 
    inputPort_4_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(14) & inputPort_4_Daemon_CP_609_elements(68);
      gj_inputPort_4_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	37 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11: 	39 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_sample_start__ps
      -- 
    inputPort_4_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(9) & inputPort_4_Daemon_CP_609_elements(15) & inputPort_4_Daemon_CP_609_elements(37) & inputPort_4_Daemon_CP_609_elements(14);
      gj_inputPort_4_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	40 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	69 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	37 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_346_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_sample_completed_
      -- 
    inputPort_4_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(17) & inputPort_4_Daemon_CP_609_elements(35) & inputPort_4_Daemon_CP_609_elements(40);
      gj_inputPort_4_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	32 
    -- CP-element group 13: 	38 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13: 	41 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/aggregated_phi_update_req
      -- 
    inputPort_4_Daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(16) & inputPort_4_Daemon_CP_609_elements(32) & inputPort_4_Daemon_CP_609_elements(38);
      gj_inputPort_4_Daemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	36 
    -- CP-element group 14: 	42 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/aggregated_phi_update_ack
      -- 
    inputPort_4_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(18) & inputPort_4_Daemon_CP_609_elements(36) & inputPort_4_Daemon_CP_609_elements(42);
      gj_inputPort_4_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_sample_start_
      -- 
    inputPort_4_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(9) & inputPort_4_Daemon_CP_609_elements(12);
      gj_inputPort_4_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	57 
    -- CP-element group 16: 	60 
    -- CP-element group 16: 	63 
    -- CP-element group 16: 	66 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_update_start_
      -- 
    inputPort_4_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(9) & inputPort_4_Daemon_CP_609_elements(57) & inputPort_4_Daemon_CP_609_elements(60) & inputPort_4_Daemon_CP_609_elements(63) & inputPort_4_Daemon_CP_609_elements(66);
      gj_inputPort_4_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_sample_completed__ps
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	56 
    -- CP-element group 18: 	59 
    -- CP-element group 18: 	62 
    -- CP-element group 18: 	65 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_update_completed_
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_loopback_trigger
      -- 
    inputPort_4_Daemon_CP_609_elements(19) <= inputPort_4_Daemon_CP_609_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_loopback_sample_req_ps
      -- 
    phi_stmt_341_loopback_sample_req_648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_341_loopback_sample_req_648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(20), ack => phi_stmt_341_req_1); -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_entry_trigger
      -- 
    inputPort_4_Daemon_CP_609_elements(21) <= inputPort_4_Daemon_CP_609_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_entry_sample_req_ps
      -- 
    phi_stmt_341_entry_sample_req_651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_341_entry_sample_req_651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(22), ack => phi_stmt_341_req_0); -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_phi_mux_ack_ps
      -- 
    phi_stmt_341_phi_mux_ack_654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_341_ack_0, ack => inputPort_4_Daemon_CP_609_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/type_cast_344_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/type_cast_344_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/type_cast_344_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/type_cast_344_sample_completed_
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/type_cast_344_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/type_cast_344_update_start_
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/type_cast_344_update_completed__ps
      -- 
    inputPort_4_Daemon_CP_609_elements(26) <= inputPort_4_Daemon_CP_609_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/type_cast_344_update_completed_
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => inputPort_4_Daemon_CP_609_elements(25), ack => inputPort_4_Daemon_CP_609_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_Sample/req
      -- 
    req_675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(28), ack => next_count_down_376_345_buf_req_0); -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_update_start_
      -- CP-element group 29: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_Update/req
      -- 
    req_680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(29), ack => next_count_down_376_345_buf_req_1); -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_Sample/ack
      -- 
    ack_676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_376_345_buf_ack_0, ack => inputPort_4_Daemon_CP_609_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_Update/ack
      -- 
    ack_681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_376_345_buf_ack_1, ack => inputPort_4_Daemon_CP_609_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	57 
    -- CP-element group 32: 	60 
    -- CP-element group 32: 	63 
    -- CP-element group 32: 	66 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_346_update_start_
      -- 
    inputPort_4_Daemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(9) & inputPort_4_Daemon_CP_609_elements(57) & inputPort_4_Daemon_CP_609_elements(60) & inputPort_4_Daemon_CP_609_elements(63) & inputPort_4_Daemon_CP_609_elements(66);
      gj_inputPort_4_Daemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/RPIPE_in_data_4_348_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/RPIPE_in_data_4_348_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/RPIPE_in_data_4_348_Sample/rr
      -- 
    rr_694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(33), ack => RPIPE_in_data_4_348_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(11) & inputPort_4_Daemon_CP_609_elements(36);
      gj_inputPort_4_Daemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	13 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/RPIPE_in_data_4_348_update_start_
      -- CP-element group 34: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/RPIPE_in_data_4_348_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/RPIPE_in_data_4_348_Update/cr
      -- 
    cr_699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(34), ack => RPIPE_in_data_4_348_inst_req_1); -- 
    inputPort_4_Daemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(13) & inputPort_4_Daemon_CP_609_elements(35);
      gj_inputPort_4_Daemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/RPIPE_in_data_4_348_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/RPIPE_in_data_4_348_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/RPIPE_in_data_4_348_Sample/ra
      -- 
    ra_695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_4_348_inst_ack_0, ack => inputPort_4_Daemon_CP_609_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	56 
    -- CP-element group 36: 	59 
    -- CP-element group 36: 	62 
    -- CP-element group 36: 	65 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_346_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/RPIPE_in_data_4_348_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/RPIPE_in_data_4_348_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/RPIPE_in_data_4_348_Update/ca
      -- 
    ca_700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_4_348_inst_ack_1, ack => inputPort_4_Daemon_CP_609_elements(36)); -- 
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	9 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	12 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	11 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_sample_start_
      -- 
    inputPort_4_Daemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(9) & inputPort_4_Daemon_CP_609_elements(12);
      gj_inputPort_4_Daemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	9 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	57 
    -- CP-element group 38: 	60 
    -- CP-element group 38: 	63 
    -- CP-element group 38: 	66 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	13 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_update_start_
      -- 
    inputPort_4_Daemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(9) & inputPort_4_Daemon_CP_609_elements(57) & inputPort_4_Daemon_CP_609_elements(60) & inputPort_4_Daemon_CP_609_elements(63) & inputPort_4_Daemon_CP_609_elements(66);
      gj_inputPort_4_Daemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	11 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_sample_start__ps
      -- 
    inputPort_4_Daemon_CP_609_elements(39) <= inputPort_4_Daemon_CP_609_elements(11);
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	12 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_sample_completed__ps
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	13 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_update_start__ps
      -- 
    inputPort_4_Daemon_CP_609_elements(41) <= inputPort_4_Daemon_CP_609_elements(13);
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	14 
    -- CP-element group 42: 	56 
    -- CP-element group 42: 	59 
    -- CP-element group 42: 	62 
    -- CP-element group 42: 	65 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_update_completed__ps
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	7 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_loopback_trigger
      -- 
    inputPort_4_Daemon_CP_609_elements(43) <= inputPort_4_Daemon_CP_609_elements(7);
    -- CP-element group 44:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_loopback_sample_req
      -- CP-element group 44: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_loopback_sample_req_ps
      -- 
    phi_stmt_349_loopback_sample_req_710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_349_loopback_sample_req_710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(44), ack => phi_stmt_349_req_1); -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	8 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_entry_trigger
      -- 
    inputPort_4_Daemon_CP_609_elements(45) <= inputPort_4_Daemon_CP_609_elements(8);
    -- CP-element group 46:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_entry_sample_req
      -- CP-element group 46: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_entry_sample_req_ps
      -- 
    phi_stmt_349_entry_sample_req_713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_349_entry_sample_req_713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(46), ack => phi_stmt_349_req_0); -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_phi_mux_ack
      -- CP-element group 47: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_phi_mux_ack_ps
      -- 
    phi_stmt_349_phi_mux_ack_716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_349_ack_0, ack => inputPort_4_Daemon_CP_609_elements(47)); -- 
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/konst_351_sample_start__ps
      -- CP-element group 48: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/konst_351_sample_completed__ps
      -- CP-element group 48: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/konst_351_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/konst_351_sample_completed_
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/konst_351_update_start__ps
      -- CP-element group 49: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/konst_351_update_start_
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/konst_351_update_completed__ps
      -- 
    inputPort_4_Daemon_CP_609_elements(50) <= inputPort_4_Daemon_CP_609_elements(51);
    -- CP-element group 51:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	50 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/konst_351_update_completed_
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(51) is a control-delay.
    cp_element_51_delay: control_delay_element  generic map(name => " 51_delay", delay_value => 1)  port map(req => inputPort_4_Daemon_CP_609_elements(49), ack => inputPort_4_Daemon_CP_609_elements(51), clk => clk, reset =>reset);
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_Sample/req
      -- 
    req_737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(52), ack => next_last_dest_id_382_352_buf_req_0); -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_update_start_
      -- CP-element group 53: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_Update/req
      -- 
    req_742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(53), ack => next_last_dest_id_382_352_buf_req_1); -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_Sample/ack
      -- 
    ack_738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_382_352_buf_ack_0, ack => inputPort_4_Daemon_CP_609_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_Update/ack
      -- 
    ack_743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_382_352_buf_ack_1, ack => inputPort_4_Daemon_CP_609_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	18 
    -- CP-element group 56: 	36 
    -- CP-element group 56: 	42 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_1_394_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_1_394_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_1_394_Sample/req
      -- 
    req_752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(56), ack => WPIPE_noblock_obuf_4_1_394_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(18) & inputPort_4_Daemon_CP_609_elements(36) & inputPort_4_Daemon_CP_609_elements(42) & inputPort_4_Daemon_CP_609_elements(58);
      gj_inputPort_4_Daemon_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	16 
    -- CP-element group 57: 	32 
    -- CP-element group 57: 	38 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_1_394_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_1_394_update_start_
      -- CP-element group 57: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_1_394_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_1_394_Sample/ack
      -- CP-element group 57: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_1_394_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_1_394_Update/req
      -- 
    ack_753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_1_394_inst_ack_0, ack => inputPort_4_Daemon_CP_609_elements(57)); -- 
    req_757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(57), ack => WPIPE_noblock_obuf_4_1_394_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	69 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_1_394_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_1_394_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_1_394_Update/ack
      -- 
    ack_758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_1_394_inst_ack_1, ack => inputPort_4_Daemon_CP_609_elements(58)); -- 
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	18 
    -- CP-element group 59: 	36 
    -- CP-element group 59: 	42 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_2_403_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_2_403_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_2_403_Sample/req
      -- 
    req_766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(59), ack => WPIPE_noblock_obuf_4_2_403_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(18) & inputPort_4_Daemon_CP_609_elements(36) & inputPort_4_Daemon_CP_609_elements(42) & inputPort_4_Daemon_CP_609_elements(61);
      gj_inputPort_4_Daemon_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	16 
    -- CP-element group 60: 	32 
    -- CP-element group 60: 	38 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_2_403_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_2_403_update_start_
      -- CP-element group 60: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_2_403_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_2_403_Sample/ack
      -- CP-element group 60: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_2_403_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_2_403_Update/req
      -- 
    ack_767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_2_403_inst_ack_0, ack => inputPort_4_Daemon_CP_609_elements(60)); -- 
    req_771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(60), ack => WPIPE_noblock_obuf_4_2_403_inst_req_1); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	69 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_2_403_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_2_403_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_2_403_Update/ack
      -- 
    ack_772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_2_403_inst_ack_1, ack => inputPort_4_Daemon_CP_609_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	18 
    -- CP-element group 62: 	36 
    -- CP-element group 62: 	42 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_3_412_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_3_412_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_3_412_Sample/req
      -- 
    req_780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(62), ack => WPIPE_noblock_obuf_4_3_412_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(18) & inputPort_4_Daemon_CP_609_elements(36) & inputPort_4_Daemon_CP_609_elements(42) & inputPort_4_Daemon_CP_609_elements(64);
      gj_inputPort_4_Daemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	16 
    -- CP-element group 63: 	32 
    -- CP-element group 63: 	38 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_3_412_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_3_412_update_start_
      -- CP-element group 63: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_3_412_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_3_412_Sample/ack
      -- CP-element group 63: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_3_412_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_3_412_Update/req
      -- 
    ack_781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_3_412_inst_ack_0, ack => inputPort_4_Daemon_CP_609_elements(63)); -- 
    req_785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(63), ack => WPIPE_noblock_obuf_4_3_412_inst_req_1); -- 
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	69 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_3_412_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_3_412_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_3_412_Update/ack
      -- 
    ack_786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_3_412_inst_ack_1, ack => inputPort_4_Daemon_CP_609_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	18 
    -- CP-element group 65: 	36 
    -- CP-element group 65: 	42 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_4_421_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_4_421_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_4_421_Sample/req
      -- 
    req_794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(65), ack => WPIPE_noblock_obuf_4_4_421_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(18) & inputPort_4_Daemon_CP_609_elements(36) & inputPort_4_Daemon_CP_609_elements(42) & inputPort_4_Daemon_CP_609_elements(67);
      gj_inputPort_4_Daemon_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	16 
    -- CP-element group 66: 	32 
    -- CP-element group 66: 	38 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_4_421_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_4_421_update_start_
      -- CP-element group 66: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_4_421_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_4_421_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_4_421_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_4_421_Update/req
      -- 
    ack_795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_4_421_inst_ack_0, ack => inputPort_4_Daemon_CP_609_elements(66)); -- 
    req_799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(66), ack => WPIPE_noblock_obuf_4_4_421_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_4_421_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_4_421_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_4_421_Update/ack
      -- 
    ack_800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_4_421_inst_ack_1, ack => inputPort_4_Daemon_CP_609_elements(67)); -- 
    -- CP-element group 68:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	9 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	10 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(68) is a control-delay.
    cp_element_68_delay: control_delay_element  generic map(name => " 68_delay", delay_value => 1)  port map(req => inputPort_4_Daemon_CP_609_elements(9), ack => inputPort_4_Daemon_CP_609_elements(68), clk => clk, reset =>reset);
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	12 
    -- CP-element group 69: 	58 
    -- CP-element group 69: 	61 
    -- CP-element group 69: 	64 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	6 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/$exit
      -- 
    inputPort_4_Daemon_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(12) & inputPort_4_Daemon_CP_609_elements(58) & inputPort_4_Daemon_CP_609_elements(61) & inputPort_4_Daemon_CP_609_elements(64) & inputPort_4_Daemon_CP_609_elements(67);
      gj_inputPort_4_Daemon_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	5 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_338/do_while_stmt_339/loop_exit/$exit
      -- CP-element group 70: 	 branch_block_stmt_338/do_while_stmt_339/loop_exit/ack
      -- 
    ack_805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_339_branch_ack_0, ack => inputPort_4_Daemon_CP_609_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	5 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_338/do_while_stmt_339/loop_taken/$exit
      -- CP-element group 71: 	 branch_block_stmt_338/do_while_stmt_339/loop_taken/ack
      -- 
    ack_809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_339_branch_ack_1, ack => inputPort_4_Daemon_CP_609_elements(71)); -- 
    -- CP-element group 72:  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	3 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	1 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_338/do_while_stmt_339/$exit
      -- 
    inputPort_4_Daemon_CP_609_elements(72) <= inputPort_4_Daemon_CP_609_elements(3);
    inputPort_4_Daemon_do_while_stmt_339_terminator_810: loop_terminator -- 
      generic map (name => " inputPort_4_Daemon_do_while_stmt_339_terminator_810", max_iterations_in_flight =>7) 
      port map(loop_body_exit => inputPort_4_Daemon_CP_609_elements(6),loop_continue => inputPort_4_Daemon_CP_609_elements(71),loop_terminate => inputPort_4_Daemon_CP_609_elements(70),loop_back => inputPort_4_Daemon_CP_609_elements(4),loop_exit => inputPort_4_Daemon_CP_609_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_341_phi_seq_682_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_4_Daemon_CP_609_elements(21);
      inputPort_4_Daemon_CP_609_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_4_Daemon_CP_609_elements(24);
      inputPort_4_Daemon_CP_609_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_4_Daemon_CP_609_elements(26);
      inputPort_4_Daemon_CP_609_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_4_Daemon_CP_609_elements(19);
      inputPort_4_Daemon_CP_609_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_4_Daemon_CP_609_elements(30);
      inputPort_4_Daemon_CP_609_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_4_Daemon_CP_609_elements(31);
      inputPort_4_Daemon_CP_609_elements(20) <= phi_mux_reqs(1);
      phi_stmt_341_phi_seq_682 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_341_phi_seq_682") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_4_Daemon_CP_609_elements(11), 
          phi_sample_ack => inputPort_4_Daemon_CP_609_elements(17), 
          phi_update_req => inputPort_4_Daemon_CP_609_elements(13), 
          phi_update_ack => inputPort_4_Daemon_CP_609_elements(18), 
          phi_mux_ack => inputPort_4_Daemon_CP_609_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_349_phi_seq_744_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_4_Daemon_CP_609_elements(45);
      inputPort_4_Daemon_CP_609_elements(48)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_4_Daemon_CP_609_elements(48);
      inputPort_4_Daemon_CP_609_elements(49)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_4_Daemon_CP_609_elements(50);
      inputPort_4_Daemon_CP_609_elements(46) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_4_Daemon_CP_609_elements(43);
      inputPort_4_Daemon_CP_609_elements(52)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_4_Daemon_CP_609_elements(54);
      inputPort_4_Daemon_CP_609_elements(53)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_4_Daemon_CP_609_elements(55);
      inputPort_4_Daemon_CP_609_elements(44) <= phi_mux_reqs(1);
      phi_stmt_349_phi_seq_744 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_349_phi_seq_744") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_4_Daemon_CP_609_elements(39), 
          phi_sample_ack => inputPort_4_Daemon_CP_609_elements(40), 
          phi_update_req => inputPort_4_Daemon_CP_609_elements(41), 
          phi_update_ack => inputPort_4_Daemon_CP_609_elements(42), 
          phi_mux_ack => inputPort_4_Daemon_CP_609_elements(47), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_634_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= inputPort_4_Daemon_CP_609_elements(7);
        preds(1)  <= inputPort_4_Daemon_CP_609_elements(8);
        entry_tmerge_634 : transition_merge -- 
          generic map(name => " entry_tmerge_634")
          port map (preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal RPIPE_in_data_4_348_wire : std_logic_vector(31 downto 0);
    signal R_ONE_1_384_wire_constant : std_logic_vector(0 downto 0);
    signal SUB_u16_u16_371_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_374_wire : std_logic_vector(15 downto 0);
    signal count_down_341 : std_logic_vector(15 downto 0);
    signal data_to_outport_387 : std_logic_vector(32 downto 0);
    signal dest_id_362 : std_logic_vector(7 downto 0);
    signal input_word_346 : std_logic_vector(31 downto 0);
    signal konst_351_wire_constant : std_logic_vector(7 downto 0);
    signal konst_356_wire_constant : std_logic_vector(15 downto 0);
    signal konst_370_wire_constant : std_logic_vector(15 downto 0);
    signal konst_373_wire_constant : std_logic_vector(15 downto 0);
    signal konst_390_wire_constant : std_logic_vector(7 downto 0);
    signal konst_399_wire_constant : std_logic_vector(7 downto 0);
    signal konst_408_wire_constant : std_logic_vector(7 downto 0);
    signal konst_417_wire_constant : std_logic_vector(7 downto 0);
    signal konst_425_wire_constant : std_logic_vector(0 downto 0);
    signal last_dest_id_349 : std_logic_vector(7 downto 0);
    signal new_packet_358 : std_logic_vector(0 downto 0);
    signal next_count_down_376 : std_logic_vector(15 downto 0);
    signal next_count_down_376_345_buffered : std_logic_vector(15 downto 0);
    signal next_last_dest_id_382 : std_logic_vector(7 downto 0);
    signal next_last_dest_id_382_352_buffered : std_logic_vector(7 downto 0);
    signal pkt_length_366 : std_logic_vector(15 downto 0);
    signal send_to_1_392 : std_logic_vector(0 downto 0);
    signal send_to_2_401 : std_logic_vector(0 downto 0);
    signal send_to_3_410 : std_logic_vector(0 downto 0);
    signal send_to_4_419 : std_logic_vector(0 downto 0);
    signal type_cast_344_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    R_ONE_1_384_wire_constant <= "1";
    konst_351_wire_constant <= "00000000";
    konst_356_wire_constant <= "0000000000000000";
    konst_370_wire_constant <= "0000000000000001";
    konst_373_wire_constant <= "0000000000000001";
    konst_390_wire_constant <= "00000001";
    konst_399_wire_constant <= "00000010";
    konst_408_wire_constant <= "00000011";
    konst_417_wire_constant <= "00000100";
    konst_425_wire_constant <= "1";
    type_cast_344_wire_constant <= "0000000000000000";
    phi_stmt_341: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_344_wire_constant & next_count_down_376_345_buffered;
      req <= phi_stmt_341_req_0 & phi_stmt_341_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_341",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_341_ack_0,
          idata => idata,
          odata => count_down_341,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_341
    phi_stmt_349: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_351_wire_constant & next_last_dest_id_382_352_buffered;
      req <= phi_stmt_349_req_0 & phi_stmt_349_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_349",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_349_ack_0,
          idata => idata,
          odata => last_dest_id_349,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_349
    -- flow-through select operator MUX_375_inst
    next_count_down_376 <= SUB_u16_u16_371_wire when (new_packet_358(0) /=  '0') else SUB_u16_u16_374_wire;
    -- flow-through select operator MUX_381_inst
    next_last_dest_id_382 <= dest_id_362 when (new_packet_358(0) /=  '0') else last_dest_id_349;
    -- flow-through slice operator slice_361_inst
    dest_id_362 <= input_word_346(31 downto 24);
    -- flow-through slice operator slice_365_inst
    pkt_length_366 <= input_word_346(23 downto 8);
    next_count_down_376_345_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_count_down_376_345_buf_req_0;
      next_count_down_376_345_buf_ack_0<= wack(0);
      rreq(0) <= next_count_down_376_345_buf_req_1;
      next_count_down_376_345_buf_ack_1<= rack(0);
      next_count_down_376_345_buf : InterlockBuffer generic map ( -- 
        name => "next_count_down_376_345_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_count_down_376,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_count_down_376_345_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_last_dest_id_382_352_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_last_dest_id_382_352_buf_req_0;
      next_last_dest_id_382_352_buf_ack_0<= wack(0);
      rreq(0) <= next_last_dest_id_382_352_buf_req_1;
      next_last_dest_id_382_352_buf_ack_1<= rack(0);
      next_last_dest_id_382_352_buf : InterlockBuffer generic map ( -- 
        name => "next_last_dest_id_382_352_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_last_dest_id_382,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_last_dest_id_382_352_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_346
    process(RPIPE_in_data_4_348_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := RPIPE_in_data_4_348_wire(31 downto 0);
      input_word_346 <= tmp_var; -- 
    end process;
    do_while_stmt_339_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_425_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_339_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_339_branch_req_0,
          ack0 => do_while_stmt_339_branch_ack_0,
          ack1 => do_while_stmt_339_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator CONCAT_u1_u33_386_inst
    process(R_ONE_1_384_wire_constant, input_word_346) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ONE_1_384_wire_constant, input_word_346, tmp_var);
      data_to_outport_387 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_357_inst
    process(count_down_341) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(count_down_341, konst_356_wire_constant, tmp_var);
      new_packet_358 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_391_inst
    process(next_last_dest_id_382) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_382, konst_390_wire_constant, tmp_var);
      send_to_1_392 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_400_inst
    process(next_last_dest_id_382) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_382, konst_399_wire_constant, tmp_var);
      send_to_2_401 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_409_inst
    process(next_last_dest_id_382) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_382, konst_408_wire_constant, tmp_var);
      send_to_3_410 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_418_inst
    process(next_last_dest_id_382) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_382, konst_417_wire_constant, tmp_var);
      send_to_4_419 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_371_inst
    process(pkt_length_366) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(pkt_length_366, konst_370_wire_constant, tmp_var);
      SUB_u16_u16_371_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_374_inst
    process(count_down_341) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(count_down_341, konst_373_wire_constant, tmp_var);
      SUB_u16_u16_374_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_in_data_4_348_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_in_data_4_348_inst_req_0;
      RPIPE_in_data_4_348_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_in_data_4_348_inst_req_1;
      RPIPE_in_data_4_348_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_in_data_4_348_wire <= data_out(31 downto 0);
      in_data_4_read_0_gI: SplitGuardInterface generic map(name => "in_data_4_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      in_data_4_read_0: InputPortRevised -- 
        generic map ( name => "in_data_4_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => in_data_4_pipe_read_req(0),
          oack => in_data_4_pipe_read_ack(0),
          odata => in_data_4_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_noblock_obuf_4_1_394_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_4_1_394_inst_req_0;
      WPIPE_noblock_obuf_4_1_394_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_4_1_394_inst_req_1;
      WPIPE_noblock_obuf_4_1_394_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_1_392(0);
      data_in <= data_to_outport_387;
      noblock_obuf_4_1_write_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_1_write_0: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_4_1", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_4_1_pipe_write_req(0),
          oack => noblock_obuf_4_1_pipe_write_ack(0),
          odata => noblock_obuf_4_1_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_noblock_obuf_4_2_403_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_4_2_403_inst_req_0;
      WPIPE_noblock_obuf_4_2_403_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_4_2_403_inst_req_1;
      WPIPE_noblock_obuf_4_2_403_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_2_401(0);
      data_in <= data_to_outport_387;
      noblock_obuf_4_2_write_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_2_write_1: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_4_2", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_4_2_pipe_write_req(0),
          oack => noblock_obuf_4_2_pipe_write_ack(0),
          odata => noblock_obuf_4_2_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_noblock_obuf_4_3_412_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_4_3_412_inst_req_0;
      WPIPE_noblock_obuf_4_3_412_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_4_3_412_inst_req_1;
      WPIPE_noblock_obuf_4_3_412_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_3_410(0);
      data_in <= data_to_outport_387;
      noblock_obuf_4_3_write_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_3_write_2: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_4_3", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_4_3_pipe_write_req(0),
          oack => noblock_obuf_4_3_pipe_write_ack(0),
          odata => noblock_obuf_4_3_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_noblock_obuf_4_4_421_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_4_4_421_inst_req_0;
      WPIPE_noblock_obuf_4_4_421_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_4_4_421_inst_req_1;
      WPIPE_noblock_obuf_4_4_421_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_4_419(0);
      data_in <= data_to_outport_387;
      noblock_obuf_4_4_write_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_4_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_4_write_3: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_4_4", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_4_4_pipe_write_req(0),
          oack => noblock_obuf_4_4_pipe_write_ack(0),
          odata => noblock_obuf_4_4_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end inputPort_4_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity outputPort_1_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    noblock_obuf_4_1_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_1_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_2_1_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_1_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_1_1_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_1_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_3_1_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_1_pipe_read_data : in   std_logic_vector(32 downto 0);
    out_data_1_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_1_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity outputPort_1_Daemon;
architecture outputPort_1_Daemon_arch of outputPort_1_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal outputPort_1_Daemon_CP_814_start: Boolean;
  signal outputPort_1_Daemon_CP_814_symbol: Boolean;
  -- volatile/operator module components. 
  component prioritySelect_Volatile is -- 
    port ( -- 
      down_counter : in  std_logic_vector(7 downto 0);
      active_packet : in  std_logic_vector(2 downto 0);
      pkt_priority : in  std_logic_vector(2 downto 0);
      p1_valid : in  std_logic_vector(0 downto 0);
      p2_valid : in  std_logic_vector(0 downto 0);
      p3_valid : in  std_logic_vector(0 downto 0);
      p4_valid : in  std_logic_vector(0 downto 0);
      next_active_packet : out  std_logic_vector(2 downto 0);
      next_pkt_priority : out  std_logic_vector(2 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal phi_stmt_589_ack_0 : boolean;
  signal do_while_stmt_587_branch_ack_1 : boolean;
  signal phi_stmt_593_req_1 : boolean;
  signal WPIPE_out_data_1_807_inst_req_1 : boolean;
  signal next_down_counter_700_592_buf_req_0 : boolean;
  signal WPIPE_out_data_1_807_inst_req_0 : boolean;
  signal next_down_counter_700_592_buf_ack_0 : boolean;
  signal do_while_stmt_587_branch_req_0 : boolean;
  signal do_while_stmt_587_branch_ack_0 : boolean;
  signal phi_stmt_593_req_0 : boolean;
  signal WPIPE_out_data_1_807_inst_ack_0 : boolean;
  signal phi_stmt_589_req_0 : boolean;
  signal RPIPE_noblock_obuf_1_1_597_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_1_597_inst_ack_1 : boolean;
  signal RPIPE_noblock_obuf_1_1_597_inst_req_0 : boolean;
  signal phi_stmt_598_req_1 : boolean;
  signal RPIPE_noblock_obuf_1_1_597_inst_req_1 : boolean;
  signal phi_stmt_589_req_1 : boolean;
  signal WPIPE_out_data_1_807_inst_ack_1 : boolean;
  signal next_down_counter_700_592_buf_ack_1 : boolean;
  signal next_down_counter_700_592_buf_req_1 : boolean;
  signal phi_stmt_593_ack_0 : boolean;
  signal phi_stmt_598_req_0 : boolean;
  signal phi_stmt_598_ack_0 : boolean;
  signal RPIPE_noblock_obuf_2_1_602_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_2_1_602_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_2_1_602_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_2_1_602_inst_ack_1 : boolean;
  signal phi_stmt_603_req_1 : boolean;
  signal phi_stmt_603_req_0 : boolean;
  signal phi_stmt_603_ack_0 : boolean;
  signal RPIPE_noblock_obuf_3_1_607_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_3_1_607_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_3_1_607_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_3_1_607_inst_ack_1 : boolean;
  signal phi_stmt_608_req_1 : boolean;
  signal phi_stmt_608_req_0 : boolean;
  signal phi_stmt_608_ack_0 : boolean;
  signal RPIPE_noblock_obuf_4_1_612_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_4_1_612_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_4_1_612_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_4_1_612_inst_ack_1 : boolean;
  signal phi_stmt_613_req_1 : boolean;
  signal phi_stmt_613_req_0 : boolean;
  signal phi_stmt_613_ack_0 : boolean;
  signal next_active_packet_680_616_buf_req_0 : boolean;
  signal next_active_packet_680_616_buf_ack_0 : boolean;
  signal next_active_packet_680_616_buf_req_1 : boolean;
  signal next_active_packet_680_616_buf_ack_1 : boolean;
  signal phi_stmt_617_req_1 : boolean;
  signal phi_stmt_617_req_0 : boolean;
  signal phi_stmt_617_ack_0 : boolean;
  signal next_pkt_priority_680_620_buf_req_0 : boolean;
  signal next_pkt_priority_680_620_buf_ack_0 : boolean;
  signal next_pkt_priority_680_620_buf_req_1 : boolean;
  signal next_pkt_priority_680_620_buf_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "outputPort_1_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  outputPort_1_Daemon_CP_814_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "outputPort_1_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_1_Daemon_CP_814_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= outputPort_1_Daemon_CP_814_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_1_Daemon_CP_814_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  outputPort_1_Daemon_CP_814: Block -- control-path 
    signal outputPort_1_Daemon_CP_814_elements: BooleanArray(161 downto 0);
    -- 
  begin -- 
    outputPort_1_Daemon_CP_814_elements(0) <= outputPort_1_Daemon_CP_814_start;
    outputPort_1_Daemon_CP_814_symbol <= outputPort_1_Daemon_CP_814_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_586/branch_block_stmt_586__entry__
      -- CP-element group 0: 	 branch_block_stmt_586/do_while_stmt_587__entry__
      -- CP-element group 0: 	 branch_block_stmt_586/$entry
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	161 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_586/branch_block_stmt_586__exit__
      -- CP-element group 1: 	 branch_block_stmt_586/do_while_stmt_587__exit__
      -- CP-element group 1: 	 branch_block_stmt_586/$exit
      -- CP-element group 1: 	 $exit
      -- 
    outputPort_1_Daemon_CP_814_elements(1) <= outputPort_1_Daemon_CP_814_elements(161);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587__entry__
      -- CP-element group 2: 	 branch_block_stmt_586/do_while_stmt_587/$entry
      -- 
    outputPort_1_Daemon_CP_814_elements(2) <= outputPort_1_Daemon_CP_814_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	161 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587__exit__
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_586/do_while_stmt_587/loop_back
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	160 
    -- CP-element group 5: 	159 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_586/do_while_stmt_587/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_586/do_while_stmt_587/condition_done
      -- CP-element group 5: 	 branch_block_stmt_586/do_while_stmt_587/loop_taken/$entry
      -- 
    outputPort_1_Daemon_CP_814_elements(5) <= outputPort_1_Daemon_CP_814_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	158 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_586/do_while_stmt_587/loop_body_done
      -- 
    outputPort_1_Daemon_CP_814_elements(6) <= outputPort_1_Daemon_CP_814_elements(158);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	38 
    -- CP-element group 7: 	59 
    -- CP-element group 7: 	80 
    -- CP-element group 7: 	101 
    -- CP-element group 7: 	122 
    -- CP-element group 7: 	141 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/back_edge_to_loop_body
      -- 
    outputPort_1_Daemon_CP_814_elements(7) <= outputPort_1_Daemon_CP_814_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	40 
    -- CP-element group 8: 	61 
    -- CP-element group 8: 	82 
    -- CP-element group 8: 	103 
    -- CP-element group 8: 	124 
    -- CP-element group 8: 	143 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/first_time_through_loop_body
      -- 
    outputPort_1_Daemon_CP_814_elements(8) <= outputPort_1_Daemon_CP_814_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	33 
    -- CP-element group 9: 	53 
    -- CP-element group 9: 	54 
    -- CP-element group 9: 	74 
    -- CP-element group 9: 	75 
    -- CP-element group 9: 	95 
    -- CP-element group 9: 	96 
    -- CP-element group 9: 	116 
    -- CP-element group 9: 	117 
    -- CP-element group 9: 	135 
    -- CP-element group 9: 	136 
    -- CP-element group 9: 	157 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/loop_body_start
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	157 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/condition_evaluated
      -- 
    condition_evaluated_838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(10), ack => do_while_stmt_587_branch_req_0); -- 
    outputPort_1_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(14) & outputPort_1_Daemon_CP_814_elements(157);
      gj_outputPort_1_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	32 
    -- CP-element group 11: 	53 
    -- CP-element group 11: 	74 
    -- CP-element group 11: 	95 
    -- CP-element group 11: 	116 
    -- CP-element group 11: 	135 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	55 
    -- CP-element group 11: 	76 
    -- CP-element group 11: 	97 
    -- CP-element group 11: 	118 
    -- CP-element group 11: 	137 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_589_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/aggregated_phi_sample_req
      -- 
    outputPort_1_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(15) & outputPort_1_Daemon_CP_814_elements(32) & outputPort_1_Daemon_CP_814_elements(53) & outputPort_1_Daemon_CP_814_elements(74) & outputPort_1_Daemon_CP_814_elements(95) & outputPort_1_Daemon_CP_814_elements(116) & outputPort_1_Daemon_CP_814_elements(135) & outputPort_1_Daemon_CP_814_elements(14);
      gj_outputPort_1_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	56 
    -- CP-element group 12: 	77 
    -- CP-element group 12: 	98 
    -- CP-element group 12: 	119 
    -- CP-element group 12: 	138 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	158 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	32 
    -- CP-element group 12: 	53 
    -- CP-element group 12: 	74 
    -- CP-element group 12: 	95 
    -- CP-element group 12: 	116 
    -- CP-element group 12: 	135 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_598_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_593_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_589_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_603_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_608_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_613_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_617_sample_completed_
      -- 
    outputPort_1_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(17) & outputPort_1_Daemon_CP_814_elements(35) & outputPort_1_Daemon_CP_814_elements(56) & outputPort_1_Daemon_CP_814_elements(77) & outputPort_1_Daemon_CP_814_elements(98) & outputPort_1_Daemon_CP_814_elements(119) & outputPort_1_Daemon_CP_814_elements(138);
      gj_outputPort_1_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	33 
    -- CP-element group 13: 	54 
    -- CP-element group 13: 	75 
    -- CP-element group 13: 	96 
    -- CP-element group 13: 	117 
    -- CP-element group 13: 	136 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	36 
    -- CP-element group 13: 	57 
    -- CP-element group 13: 	78 
    -- CP-element group 13: 	99 
    -- CP-element group 13: 	120 
    -- CP-element group 13: 	139 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_589_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/aggregated_phi_update_req
      -- 
    outputPort_1_Daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(16) & outputPort_1_Daemon_CP_814_elements(33) & outputPort_1_Daemon_CP_814_elements(54) & outputPort_1_Daemon_CP_814_elements(75) & outputPort_1_Daemon_CP_814_elements(96) & outputPort_1_Daemon_CP_814_elements(117) & outputPort_1_Daemon_CP_814_elements(136);
      gj_outputPort_1_Daemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	37 
    -- CP-element group 14: 	58 
    -- CP-element group 14: 	79 
    -- CP-element group 14: 	100 
    -- CP-element group 14: 	121 
    -- CP-element group 14: 	140 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/aggregated_phi_update_ack
      -- 
    outputPort_1_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(18) & outputPort_1_Daemon_CP_814_elements(37) & outputPort_1_Daemon_CP_814_elements(58) & outputPort_1_Daemon_CP_814_elements(79) & outputPort_1_Daemon_CP_814_elements(100) & outputPort_1_Daemon_CP_814_elements(121) & outputPort_1_Daemon_CP_814_elements(140);
      gj_outputPort_1_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_589_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	155 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_589_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(155);
      gj_outputPort_1_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_589_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	154 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_589_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_589_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_589_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(19) <= outputPort_1_Daemon_CP_814_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_589_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_589_loopback_sample_req_ps
      -- 
    phi_stmt_589_loopback_sample_req_853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_589_loopback_sample_req_853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(20), ack => phi_stmt_589_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_589_entry_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(21) <= outputPort_1_Daemon_CP_814_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_589_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_589_entry_sample_req_ps
      -- 
    phi_stmt_589_entry_sample_req_856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_589_entry_sample_req_856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(22), ack => phi_stmt_589_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_589_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_589_phi_mux_ack_ps
      -- 
    phi_stmt_589_phi_mux_ack_859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_589_ack_0, ack => outputPort_1_Daemon_CP_814_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_8_591_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_8_591_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_8_591_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_8_591_sample_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_8_591_update_start_
      -- CP-element group 25: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_8_591_update_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_8_591_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(26) <= outputPort_1_Daemon_CP_814_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_8_591_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_814_elements(25), ack => outputPort_1_Daemon_CP_814_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_down_counter_592_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_down_counter_592_Sample/req
      -- CP-element group 28: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_down_counter_592_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_down_counter_592_sample_start__ps
      -- 
    req_880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(28), ack => next_down_counter_700_592_buf_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_down_counter_592_update_start_
      -- CP-element group 29: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_down_counter_592_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_down_counter_592_Update/req
      -- CP-element group 29: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_down_counter_592_Update/$entry
      -- 
    req_885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(29), ack => next_down_counter_700_592_buf_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_down_counter_592_Sample/ack
      -- CP-element group 30: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_down_counter_592_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_down_counter_592_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_down_counter_592_sample_completed__ps
      -- 
    ack_881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_700_592_buf_ack_0, ack => outputPort_1_Daemon_CP_814_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_down_counter_592_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_down_counter_592_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_down_counter_592_Update/ack
      -- CP-element group 31: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_down_counter_592_Update/$exit
      -- 
    ack_886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_700_592_buf_ack_1, ack => outputPort_1_Daemon_CP_814_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	12 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	11 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_593_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	9 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	155 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	13 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_593_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(155);
      gj_outputPort_1_Daemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	11 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_593_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(34) <= outputPort_1_Daemon_CP_814_elements(11);
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_593_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(35) is bound as output of CP function.
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	13 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_593_update_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(36) <= outputPort_1_Daemon_CP_814_elements(13);
    -- CP-element group 37:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	14 
    -- CP-element group 37: 	154 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_593_update_completed__ps
      -- CP-element group 37: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_593_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	7 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_593_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(38) <= outputPort_1_Daemon_CP_814_elements(7);
    -- CP-element group 39:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_593_loopback_sample_req
      -- CP-element group 39: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_593_loopback_sample_req_ps
      -- 
    phi_stmt_593_loopback_sample_req_897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_593_loopback_sample_req_897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(39), ack => phi_stmt_593_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	8 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_593_entry_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(40) <= outputPort_1_Daemon_CP_814_elements(8);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_593_entry_sample_req
      -- CP-element group 41: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_593_entry_sample_req_ps
      -- 
    phi_stmt_593_entry_sample_req_900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_593_entry_sample_req_900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(41), ack => phi_stmt_593_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(41) is bound as output of CP function.
    -- CP-element group 42:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_593_phi_mux_ack_ps
      -- CP-element group 42: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_593_phi_mux_ack
      -- 
    phi_stmt_593_phi_mux_ack_903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_593_ack_0, ack => outputPort_1_Daemon_CP_814_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (4) 
      -- CP-element group 43: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_595_sample_completed__ps
      -- CP-element group 43: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_595_sample_start__ps
      -- CP-element group 43: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_595_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_595_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_595_update_start__ps
      -- CP-element group 44: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_595_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(44) is bound as output of CP function.
    -- CP-element group 45:  join  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_595_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(45) <= outputPort_1_Daemon_CP_814_elements(46);
    -- CP-element group 46:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	45 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_595_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(46) is a control-delay.
    cp_element_46_delay: control_delay_element  generic map(name => " 46_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_814_elements(44), ack => outputPort_1_Daemon_CP_814_elements(46), clk => clk, reset =>reset);
    -- CP-element group 47:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_1_1_597_sample_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_1_1_597_update_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: marked-predecessors 
    -- CP-element group 49: 	52 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_1_1_597_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_1_1_597_Sample/rr
      -- CP-element group 49: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_1_1_597_sample_start_
      -- 
    rr_924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(49), ack => RPIPE_noblock_obuf_1_1_597_inst_req_0); -- 
    outputPort_1_Daemon_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(47) & outputPort_1_Daemon_CP_814_elements(52);
      gj_outputPort_1_Daemon_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: 	51 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_1_1_597_update_start_
      -- CP-element group 50: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_1_1_597_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_1_1_597_Update/cr
      -- 
    cr_929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(50), ack => RPIPE_noblock_obuf_1_1_597_inst_req_1); -- 
    outputPort_1_Daemon_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(48) & outputPort_1_Daemon_CP_814_elements(51);
      gj_outputPort_1_Daemon_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	50 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_1_1_597_sample_completed__ps
      -- CP-element group 51: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_1_1_597_Sample/ra
      -- CP-element group 51: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_1_1_597_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_1_1_597_sample_completed_
      -- 
    ra_925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_1_597_inst_ack_0, ack => outputPort_1_Daemon_CP_814_elements(51)); -- 
    -- CP-element group 52:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: marked-successors 
    -- CP-element group 52: 	49 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_1_1_597_update_completed__ps
      -- CP-element group 52: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_1_1_597_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_1_1_597_Update/ca
      -- CP-element group 52: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_1_1_597_Update/$exit
      -- 
    ca_930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_1_597_inst_ack_1, ack => outputPort_1_Daemon_CP_814_elements(52)); -- 
    -- CP-element group 53:  join  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	9 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	12 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	11 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_598_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	9 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	155 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	13 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_598_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(155);
      gj_outputPort_1_Daemon_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	11 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_598_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(55) <= outputPort_1_Daemon_CP_814_elements(11);
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	12 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_598_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(56) is bound as output of CP function.
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	13 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_598_update_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(57) <= outputPort_1_Daemon_CP_814_elements(13);
    -- CP-element group 58:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	14 
    -- CP-element group 58: 	154 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_598_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_598_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	7 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_598_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(59) <= outputPort_1_Daemon_CP_814_elements(7);
    -- CP-element group 60:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_598_loopback_sample_req
      -- CP-element group 60: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_598_loopback_sample_req_ps
      -- 
    phi_stmt_598_loopback_sample_req_941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_598_loopback_sample_req_941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(60), ack => phi_stmt_598_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	8 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_598_entry_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(61) <= outputPort_1_Daemon_CP_814_elements(8);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_598_entry_sample_req
      -- CP-element group 62: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_598_entry_sample_req_ps
      -- 
    phi_stmt_598_entry_sample_req_944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_598_entry_sample_req_944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(62), ack => phi_stmt_598_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_598_phi_mux_ack
      -- CP-element group 63: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_598_phi_mux_ack_ps
      -- 
    phi_stmt_598_phi_mux_ack_947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_598_ack_0, ack => outputPort_1_Daemon_CP_814_elements(63)); -- 
    -- CP-element group 64:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (4) 
      -- CP-element group 64: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_600_sample_start__ps
      -- CP-element group 64: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_600_sample_completed__ps
      -- CP-element group 64: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_600_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_600_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_600_update_start__ps
      -- CP-element group 65: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_600_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(65) is bound as output of CP function.
    -- CP-element group 66:  join  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_600_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(66) <= outputPort_1_Daemon_CP_814_elements(67);
    -- CP-element group 67:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	66 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_600_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(67) is a control-delay.
    cp_element_67_delay: control_delay_element  generic map(name => " 67_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_814_elements(65), ack => outputPort_1_Daemon_CP_814_elements(67), clk => clk, reset =>reset);
    -- CP-element group 68:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_2_1_602_sample_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_2_1_602_update_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(69) is bound as output of CP function.
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	73 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_2_1_602_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_2_1_602_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_2_1_602_Sample/rr
      -- 
    rr_968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(70), ack => RPIPE_noblock_obuf_2_1_602_inst_req_0); -- 
    outputPort_1_Daemon_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(68) & outputPort_1_Daemon_CP_814_elements(73);
      gj_outputPort_1_Daemon_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: 	72 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_2_1_602_update_start_
      -- CP-element group 71: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_2_1_602_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_2_1_602_Update/cr
      -- 
    cr_973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(71), ack => RPIPE_noblock_obuf_2_1_602_inst_req_1); -- 
    outputPort_1_Daemon_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(69) & outputPort_1_Daemon_CP_814_elements(72);
      gj_outputPort_1_Daemon_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	71 
    -- CP-element group 72:  members (4) 
      -- CP-element group 72: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_2_1_602_sample_completed__ps
      -- CP-element group 72: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_2_1_602_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_2_1_602_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_2_1_602_Sample/ra
      -- 
    ra_969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_1_602_inst_ack_0, ack => outputPort_1_Daemon_CP_814_elements(72)); -- 
    -- CP-element group 73:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: marked-successors 
    -- CP-element group 73: 	70 
    -- CP-element group 73:  members (4) 
      -- CP-element group 73: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_2_1_602_update_completed__ps
      -- CP-element group 73: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_2_1_602_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_2_1_602_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_2_1_602_Update/ca
      -- 
    ca_974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_1_602_inst_ack_1, ack => outputPort_1_Daemon_CP_814_elements(73)); -- 
    -- CP-element group 74:  join  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	9 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	12 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	11 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_603_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	9 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	155 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	13 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_603_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(155);
      gj_outputPort_1_Daemon_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	11 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_603_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(76) <= outputPort_1_Daemon_CP_814_elements(11);
    -- CP-element group 77:  join  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	12 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_603_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(77) is bound as output of CP function.
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	13 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_603_update_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(78) <= outputPort_1_Daemon_CP_814_elements(13);
    -- CP-element group 79:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	14 
    -- CP-element group 79: 	154 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_603_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_603_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	7 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_603_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(80) <= outputPort_1_Daemon_CP_814_elements(7);
    -- CP-element group 81:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_603_loopback_sample_req
      -- CP-element group 81: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_603_loopback_sample_req_ps
      -- 
    phi_stmt_603_loopback_sample_req_985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_603_loopback_sample_req_985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(81), ack => phi_stmt_603_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	8 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_603_entry_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(82) <= outputPort_1_Daemon_CP_814_elements(8);
    -- CP-element group 83:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_603_entry_sample_req
      -- CP-element group 83: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_603_entry_sample_req_ps
      -- 
    phi_stmt_603_entry_sample_req_988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_603_entry_sample_req_988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(83), ack => phi_stmt_603_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(83) is bound as output of CP function.
    -- CP-element group 84:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_603_phi_mux_ack_ps
      -- CP-element group 84: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_603_phi_mux_ack
      -- 
    phi_stmt_603_phi_mux_ack_991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_603_ack_0, ack => outputPort_1_Daemon_CP_814_elements(84)); -- 
    -- CP-element group 85:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (4) 
      -- CP-element group 85: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_605_sample_start__ps
      -- CP-element group 85: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_605_sample_completed__ps
      -- CP-element group 85: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_605_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_605_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_605_update_start__ps
      -- CP-element group 86: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_605_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(86) is bound as output of CP function.
    -- CP-element group 87:  join  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_605_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(87) <= outputPort_1_Daemon_CP_814_elements(88);
    -- CP-element group 88:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	87 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_605_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(88) is a control-delay.
    cp_element_88_delay: control_delay_element  generic map(name => " 88_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_814_elements(86), ack => outputPort_1_Daemon_CP_814_elements(88), clk => clk, reset =>reset);
    -- CP-element group 89:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_3_1_607_sample_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(89) is bound as output of CP function.
    -- CP-element group 90:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_3_1_607_update_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(90) is bound as output of CP function.
    -- CP-element group 91:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: marked-predecessors 
    -- CP-element group 91: 	94 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_3_1_607_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_3_1_607_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_3_1_607_Sample/rr
      -- 
    rr_1012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(91), ack => RPIPE_noblock_obuf_3_1_607_inst_req_0); -- 
    outputPort_1_Daemon_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(89) & outputPort_1_Daemon_CP_814_elements(94);
      gj_outputPort_1_Daemon_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	93 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_3_1_607_update_start_
      -- CP-element group 92: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_3_1_607_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_3_1_607_Update/cr
      -- 
    cr_1017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(92), ack => RPIPE_noblock_obuf_3_1_607_inst_req_1); -- 
    outputPort_1_Daemon_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(90) & outputPort_1_Daemon_CP_814_elements(93);
      gj_outputPort_1_Daemon_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	92 
    -- CP-element group 93:  members (4) 
      -- CP-element group 93: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_3_1_607_sample_completed__ps
      -- CP-element group 93: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_3_1_607_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_3_1_607_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_3_1_607_Sample/ra
      -- 
    ra_1013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_1_607_inst_ack_0, ack => outputPort_1_Daemon_CP_814_elements(93)); -- 
    -- CP-element group 94:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: successors 
    -- CP-element group 94: marked-successors 
    -- CP-element group 94: 	91 
    -- CP-element group 94:  members (4) 
      -- CP-element group 94: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_3_1_607_update_completed__ps
      -- CP-element group 94: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_3_1_607_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_3_1_607_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_3_1_607_Update/ca
      -- 
    ca_1018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_1_607_inst_ack_1, ack => outputPort_1_Daemon_CP_814_elements(94)); -- 
    -- CP-element group 95:  join  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	9 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	12 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	11 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_608_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	9 
    -- CP-element group 96: marked-predecessors 
    -- CP-element group 96: 	155 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	13 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_608_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(155);
      gj_outputPort_1_Daemon_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	11 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_608_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(97) <= outputPort_1_Daemon_CP_814_elements(11);
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	12 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_608_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(98) is bound as output of CP function.
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	13 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_608_update_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(99) <= outputPort_1_Daemon_CP_814_elements(13);
    -- CP-element group 100:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	14 
    -- CP-element group 100: 	154 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_608_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_608_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(100) is bound as output of CP function.
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	7 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_608_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(101) <= outputPort_1_Daemon_CP_814_elements(7);
    -- CP-element group 102:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_608_loopback_sample_req
      -- CP-element group 102: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_608_loopback_sample_req_ps
      -- 
    phi_stmt_608_loopback_sample_req_1029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_608_loopback_sample_req_1029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(102), ack => phi_stmt_608_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(102) is bound as output of CP function.
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	8 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_608_entry_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(103) <= outputPort_1_Daemon_CP_814_elements(8);
    -- CP-element group 104:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_608_entry_sample_req
      -- CP-element group 104: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_608_entry_sample_req_ps
      -- 
    phi_stmt_608_entry_sample_req_1032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_608_entry_sample_req_1032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(104), ack => phi_stmt_608_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(104) is bound as output of CP function.
    -- CP-element group 105:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_608_phi_mux_ack
      -- CP-element group 105: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_608_phi_mux_ack_ps
      -- 
    phi_stmt_608_phi_mux_ack_1035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_608_ack_0, ack => outputPort_1_Daemon_CP_814_elements(105)); -- 
    -- CP-element group 106:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (4) 
      -- CP-element group 106: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_610_sample_start__ps
      -- CP-element group 106: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_610_sample_completed__ps
      -- CP-element group 106: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_610_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_610_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_610_update_start__ps
      -- CP-element group 107: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_610_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(107) is bound as output of CP function.
    -- CP-element group 108:  join  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	109 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_610_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(108) <= outputPort_1_Daemon_CP_814_elements(109);
    -- CP-element group 109:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	108 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_33_610_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(109) is a control-delay.
    cp_element_109_delay: control_delay_element  generic map(name => " 109_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_814_elements(107), ack => outputPort_1_Daemon_CP_814_elements(109), clk => clk, reset =>reset);
    -- CP-element group 110:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_4_1_612_sample_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(110) is bound as output of CP function.
    -- CP-element group 111:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_4_1_612_update_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(111) is bound as output of CP function.
    -- CP-element group 112:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	115 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_4_1_612_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_4_1_612_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_4_1_612_Sample/rr
      -- 
    rr_1056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(112), ack => RPIPE_noblock_obuf_4_1_612_inst_req_0); -- 
    outputPort_1_Daemon_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(110) & outputPort_1_Daemon_CP_814_elements(115);
      gj_outputPort_1_Daemon_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: 	114 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_4_1_612_update_start_
      -- CP-element group 113: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_4_1_612_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_4_1_612_Update/cr
      -- 
    cr_1061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(113), ack => RPIPE_noblock_obuf_4_1_612_inst_req_1); -- 
    outputPort_1_Daemon_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(111) & outputPort_1_Daemon_CP_814_elements(114);
      gj_outputPort_1_Daemon_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	113 
    -- CP-element group 114:  members (4) 
      -- CP-element group 114: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_4_1_612_sample_completed__ps
      -- CP-element group 114: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_4_1_612_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_4_1_612_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_4_1_612_Sample/ra
      -- 
    ra_1057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_1_612_inst_ack_0, ack => outputPort_1_Daemon_CP_814_elements(114)); -- 
    -- CP-element group 115:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	112 
    -- CP-element group 115:  members (4) 
      -- CP-element group 115: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_4_1_612_update_completed__ps
      -- CP-element group 115: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_4_1_612_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_4_1_612_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/RPIPE_noblock_obuf_4_1_612_Update/ca
      -- 
    ca_1062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_1_612_inst_ack_1, ack => outputPort_1_Daemon_CP_814_elements(115)); -- 
    -- CP-element group 116:  join  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	9 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	12 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	11 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_613_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  transition  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	9 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	155 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	13 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_613_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(155);
      gj_outputPort_1_Daemon_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	11 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_613_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(118) <= outputPort_1_Daemon_CP_814_elements(11);
    -- CP-element group 119:  join  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	12 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_613_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(119) is bound as output of CP function.
    -- CP-element group 120:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	13 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_613_update_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(120) <= outputPort_1_Daemon_CP_814_elements(13);
    -- CP-element group 121:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	14 
    -- CP-element group 121: 	154 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_613_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_613_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(121) is bound as output of CP function.
    -- CP-element group 122:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	7 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_613_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(122) <= outputPort_1_Daemon_CP_814_elements(7);
    -- CP-element group 123:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_613_loopback_sample_req
      -- CP-element group 123: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_613_loopback_sample_req_ps
      -- 
    phi_stmt_613_loopback_sample_req_1073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_613_loopback_sample_req_1073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(123), ack => phi_stmt_613_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(123) is bound as output of CP function.
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	8 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_613_entry_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(124) <= outputPort_1_Daemon_CP_814_elements(8);
    -- CP-element group 125:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_613_entry_sample_req
      -- CP-element group 125: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_613_entry_sample_req_ps
      -- 
    phi_stmt_613_entry_sample_req_1076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_613_entry_sample_req_1076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(125), ack => phi_stmt_613_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(125) is bound as output of CP function.
    -- CP-element group 126:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_613_phi_mux_ack
      -- CP-element group 126: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_613_phi_mux_ack_ps
      -- 
    phi_stmt_613_phi_mux_ack_1079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_613_ack_0, ack => outputPort_1_Daemon_CP_814_elements(126)); -- 
    -- CP-element group 127:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (4) 
      -- CP-element group 127: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_3_615_sample_start__ps
      -- CP-element group 127: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_3_615_sample_completed__ps
      -- CP-element group 127: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_3_615_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_3_615_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(127) is bound as output of CP function.
    -- CP-element group 128:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_3_615_update_start__ps
      -- CP-element group 128: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_3_615_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(128) is bound as output of CP function.
    -- CP-element group 129:  join  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	130 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_3_615_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(129) <= outputPort_1_Daemon_CP_814_elements(130);
    -- CP-element group 130:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	129 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ZERO_3_615_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(130) is a control-delay.
    cp_element_130_delay: control_delay_element  generic map(name => " 130_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_814_elements(128), ack => outputPort_1_Daemon_CP_814_elements(130), clk => clk, reset =>reset);
    -- CP-element group 131:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (4) 
      -- CP-element group 131: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_active_packet_616_sample_start__ps
      -- CP-element group 131: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_active_packet_616_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_active_packet_616_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_active_packet_616_Sample/req
      -- 
    req_1100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(131), ack => next_active_packet_680_616_buf_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(131) is bound as output of CP function.
    -- CP-element group 132:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (4) 
      -- CP-element group 132: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_active_packet_616_update_start__ps
      -- CP-element group 132: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_active_packet_616_update_start_
      -- CP-element group 132: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_active_packet_616_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_active_packet_616_Update/req
      -- 
    req_1105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(132), ack => next_active_packet_680_616_buf_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(132) is bound as output of CP function.
    -- CP-element group 133:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_active_packet_616_sample_completed__ps
      -- CP-element group 133: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_active_packet_616_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_active_packet_616_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_active_packet_616_Sample/ack
      -- 
    ack_1101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_680_616_buf_ack_0, ack => outputPort_1_Daemon_CP_814_elements(133)); -- 
    -- CP-element group 134:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_active_packet_616_update_completed__ps
      -- CP-element group 134: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_active_packet_616_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_active_packet_616_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_active_packet_616_Update/ack
      -- 
    ack_1106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_680_616_buf_ack_1, ack => outputPort_1_Daemon_CP_814_elements(134)); -- 
    -- CP-element group 135:  join  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	9 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	12 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	11 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_617_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	9 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	155 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	13 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_617_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(155);
      gj_outputPort_1_Daemon_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	11 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_617_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(137) <= outputPort_1_Daemon_CP_814_elements(11);
    -- CP-element group 138:  join  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	12 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_617_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(138) is bound as output of CP function.
    -- CP-element group 139:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	13 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_617_update_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(139) <= outputPort_1_Daemon_CP_814_elements(13);
    -- CP-element group 140:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	14 
    -- CP-element group 140: 	154 
    -- CP-element group 140:  members (2) 
      -- CP-element group 140: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_617_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_617_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(140) is bound as output of CP function.
    -- CP-element group 141:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	7 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_617_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(141) <= outputPort_1_Daemon_CP_814_elements(7);
    -- CP-element group 142:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_617_loopback_sample_req
      -- CP-element group 142: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_617_loopback_sample_req_ps
      -- 
    phi_stmt_617_loopback_sample_req_1117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_617_loopback_sample_req_1117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(142), ack => phi_stmt_617_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(142) is bound as output of CP function.
    -- CP-element group 143:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	8 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_617_entry_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(143) <= outputPort_1_Daemon_CP_814_elements(8);
    -- CP-element group 144:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_617_entry_sample_req
      -- CP-element group 144: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_617_entry_sample_req_ps
      -- 
    phi_stmt_617_entry_sample_req_1120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_617_entry_sample_req_1120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(144), ack => phi_stmt_617_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_617_phi_mux_ack
      -- CP-element group 145: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/phi_stmt_617_phi_mux_ack_ps
      -- 
    phi_stmt_617_phi_mux_ack_1123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_617_ack_0, ack => outputPort_1_Daemon_CP_814_elements(145)); -- 
    -- CP-element group 146:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (4) 
      -- CP-element group 146: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ONE_3_619_sample_start__ps
      -- CP-element group 146: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ONE_3_619_sample_completed__ps
      -- CP-element group 146: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ONE_3_619_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ONE_3_619_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(146) is bound as output of CP function.
    -- CP-element group 147:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (2) 
      -- CP-element group 147: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ONE_3_619_update_start__ps
      -- CP-element group 147: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ONE_3_619_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(147) is bound as output of CP function.
    -- CP-element group 148:  join  transition  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	149 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (1) 
      -- CP-element group 148: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ONE_3_619_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(148) <= outputPort_1_Daemon_CP_814_elements(149);
    -- CP-element group 149:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	148 
    -- CP-element group 149:  members (1) 
      -- CP-element group 149: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_ONE_3_619_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(149) is a control-delay.
    cp_element_149_delay: control_delay_element  generic map(name => " 149_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_814_elements(147), ack => outputPort_1_Daemon_CP_814_elements(149), clk => clk, reset =>reset);
    -- CP-element group 150:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (4) 
      -- CP-element group 150: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_pkt_priority_620_sample_start__ps
      -- CP-element group 150: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_pkt_priority_620_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_pkt_priority_620_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_pkt_priority_620_Sample/req
      -- 
    req_1144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(150), ack => next_pkt_priority_680_620_buf_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(150) is bound as output of CP function.
    -- CP-element group 151:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (4) 
      -- CP-element group 151: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_pkt_priority_620_update_start__ps
      -- CP-element group 151: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_pkt_priority_620_update_start_
      -- CP-element group 151: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_pkt_priority_620_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_pkt_priority_620_Update/req
      -- 
    req_1149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(151), ack => next_pkt_priority_680_620_buf_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(151) is bound as output of CP function.
    -- CP-element group 152:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (4) 
      -- CP-element group 152: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_pkt_priority_620_sample_completed__ps
      -- CP-element group 152: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_pkt_priority_620_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_pkt_priority_620_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_pkt_priority_620_Sample/ack
      -- 
    ack_1145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pkt_priority_680_620_buf_ack_0, ack => outputPort_1_Daemon_CP_814_elements(152)); -- 
    -- CP-element group 153:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (4) 
      -- CP-element group 153: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_pkt_priority_620_update_completed__ps
      -- CP-element group 153: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_pkt_priority_620_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_pkt_priority_620_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/R_next_pkt_priority_620_Update/ack
      -- 
    ack_1150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pkt_priority_680_620_buf_ack_1, ack => outputPort_1_Daemon_CP_814_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	18 
    -- CP-element group 154: 	37 
    -- CP-element group 154: 	58 
    -- CP-element group 154: 	79 
    -- CP-element group 154: 	100 
    -- CP-element group 154: 	121 
    -- CP-element group 154: 	140 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/WPIPE_out_data_1_807_Sample/req
      -- CP-element group 154: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/WPIPE_out_data_1_807_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/WPIPE_out_data_1_807_sample_start_
      -- 
    req_1159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(154), ack => WPIPE_out_data_1_807_inst_req_0); -- 
    outputPort_1_Daemon_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(18) & outputPort_1_Daemon_CP_814_elements(37) & outputPort_1_Daemon_CP_814_elements(58) & outputPort_1_Daemon_CP_814_elements(79) & outputPort_1_Daemon_CP_814_elements(100) & outputPort_1_Daemon_CP_814_elements(121) & outputPort_1_Daemon_CP_814_elements(140) & outputPort_1_Daemon_CP_814_elements(156);
      gj_outputPort_1_Daemon_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	16 
    -- CP-element group 155: 	33 
    -- CP-element group 155: 	54 
    -- CP-element group 155: 	75 
    -- CP-element group 155: 	96 
    -- CP-element group 155: 	117 
    -- CP-element group 155: 	136 
    -- CP-element group 155:  members (6) 
      -- CP-element group 155: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/WPIPE_out_data_1_807_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/WPIPE_out_data_1_807_Update/req
      -- CP-element group 155: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/WPIPE_out_data_1_807_Sample/ack
      -- CP-element group 155: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/WPIPE_out_data_1_807_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/WPIPE_out_data_1_807_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/WPIPE_out_data_1_807_update_start_
      -- 
    ack_1160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_1_807_inst_ack_0, ack => outputPort_1_Daemon_CP_814_elements(155)); -- 
    req_1164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(155), ack => WPIPE_out_data_1_807_inst_req_1); -- 
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	154 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/WPIPE_out_data_1_807_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/WPIPE_out_data_1_807_Update/ack
      -- CP-element group 156: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/WPIPE_out_data_1_807_update_completed_
      -- 
    ack_1165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_1_807_inst_ack_1, ack => outputPort_1_Daemon_CP_814_elements(156)); -- 
    -- CP-element group 157:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	9 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	10 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(157) is a control-delay.
    cp_element_157_delay: control_delay_element  generic map(name => " 157_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_814_elements(9), ack => outputPort_1_Daemon_CP_814_elements(157), clk => clk, reset =>reset);
    -- CP-element group 158:  join  transition  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	12 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	6 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_586/do_while_stmt_587/do_while_stmt_587_loop_body/$exit
      -- 
    outputPort_1_Daemon_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(12) & outputPort_1_Daemon_CP_814_elements(156);
      gj_outputPort_1_Daemon_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	5 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (2) 
      -- CP-element group 159: 	 branch_block_stmt_586/do_while_stmt_587/loop_exit/ack
      -- CP-element group 159: 	 branch_block_stmt_586/do_while_stmt_587/loop_exit/$exit
      -- 
    ack_1170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_587_branch_ack_0, ack => outputPort_1_Daemon_CP_814_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	5 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (2) 
      -- CP-element group 160: 	 branch_block_stmt_586/do_while_stmt_587/loop_taken/ack
      -- CP-element group 160: 	 branch_block_stmt_586/do_while_stmt_587/loop_taken/$exit
      -- 
    ack_1174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_587_branch_ack_1, ack => outputPort_1_Daemon_CP_814_elements(160)); -- 
    -- CP-element group 161:  transition  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	3 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	1 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_586/do_while_stmt_587/$exit
      -- 
    outputPort_1_Daemon_CP_814_elements(161) <= outputPort_1_Daemon_CP_814_elements(3);
    outputPort_1_Daemon_do_while_stmt_587_terminator_1175: loop_terminator -- 
      generic map (name => " outputPort_1_Daemon_do_while_stmt_587_terminator_1175", max_iterations_in_flight =>7) 
      port map(loop_body_exit => outputPort_1_Daemon_CP_814_elements(6),loop_continue => outputPort_1_Daemon_CP_814_elements(160),loop_terminate => outputPort_1_Daemon_CP_814_elements(159),loop_back => outputPort_1_Daemon_CP_814_elements(4),loop_exit => outputPort_1_Daemon_CP_814_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_589_phi_seq_887_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_814_elements(21);
      outputPort_1_Daemon_CP_814_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_814_elements(24);
      outputPort_1_Daemon_CP_814_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_814_elements(26);
      outputPort_1_Daemon_CP_814_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_814_elements(19);
      outputPort_1_Daemon_CP_814_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_814_elements(30);
      outputPort_1_Daemon_CP_814_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_814_elements(31);
      outputPort_1_Daemon_CP_814_elements(20) <= phi_mux_reqs(1);
      phi_stmt_589_phi_seq_887 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_589_phi_seq_887") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_814_elements(11), 
          phi_sample_ack => outputPort_1_Daemon_CP_814_elements(17), 
          phi_update_req => outputPort_1_Daemon_CP_814_elements(13), 
          phi_update_ack => outputPort_1_Daemon_CP_814_elements(18), 
          phi_mux_ack => outputPort_1_Daemon_CP_814_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_593_phi_seq_931_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_814_elements(40);
      outputPort_1_Daemon_CP_814_elements(43)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_814_elements(43);
      outputPort_1_Daemon_CP_814_elements(44)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_814_elements(45);
      outputPort_1_Daemon_CP_814_elements(41) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_814_elements(38);
      outputPort_1_Daemon_CP_814_elements(47)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_814_elements(51);
      outputPort_1_Daemon_CP_814_elements(48)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_814_elements(52);
      outputPort_1_Daemon_CP_814_elements(39) <= phi_mux_reqs(1);
      phi_stmt_593_phi_seq_931 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_593_phi_seq_931") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_814_elements(34), 
          phi_sample_ack => outputPort_1_Daemon_CP_814_elements(35), 
          phi_update_req => outputPort_1_Daemon_CP_814_elements(36), 
          phi_update_ack => outputPort_1_Daemon_CP_814_elements(37), 
          phi_mux_ack => outputPort_1_Daemon_CP_814_elements(42), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_598_phi_seq_975_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_814_elements(61);
      outputPort_1_Daemon_CP_814_elements(64)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_814_elements(64);
      outputPort_1_Daemon_CP_814_elements(65)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_814_elements(66);
      outputPort_1_Daemon_CP_814_elements(62) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_814_elements(59);
      outputPort_1_Daemon_CP_814_elements(68)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_814_elements(72);
      outputPort_1_Daemon_CP_814_elements(69)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_814_elements(73);
      outputPort_1_Daemon_CP_814_elements(60) <= phi_mux_reqs(1);
      phi_stmt_598_phi_seq_975 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_598_phi_seq_975") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_814_elements(55), 
          phi_sample_ack => outputPort_1_Daemon_CP_814_elements(56), 
          phi_update_req => outputPort_1_Daemon_CP_814_elements(57), 
          phi_update_ack => outputPort_1_Daemon_CP_814_elements(58), 
          phi_mux_ack => outputPort_1_Daemon_CP_814_elements(63), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_603_phi_seq_1019_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_814_elements(82);
      outputPort_1_Daemon_CP_814_elements(85)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_814_elements(85);
      outputPort_1_Daemon_CP_814_elements(86)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_814_elements(87);
      outputPort_1_Daemon_CP_814_elements(83) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_814_elements(80);
      outputPort_1_Daemon_CP_814_elements(89)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_814_elements(93);
      outputPort_1_Daemon_CP_814_elements(90)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_814_elements(94);
      outputPort_1_Daemon_CP_814_elements(81) <= phi_mux_reqs(1);
      phi_stmt_603_phi_seq_1019 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_603_phi_seq_1019") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_814_elements(76), 
          phi_sample_ack => outputPort_1_Daemon_CP_814_elements(77), 
          phi_update_req => outputPort_1_Daemon_CP_814_elements(78), 
          phi_update_ack => outputPort_1_Daemon_CP_814_elements(79), 
          phi_mux_ack => outputPort_1_Daemon_CP_814_elements(84), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_608_phi_seq_1063_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_814_elements(103);
      outputPort_1_Daemon_CP_814_elements(106)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_814_elements(106);
      outputPort_1_Daemon_CP_814_elements(107)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_814_elements(108);
      outputPort_1_Daemon_CP_814_elements(104) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_814_elements(101);
      outputPort_1_Daemon_CP_814_elements(110)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_814_elements(114);
      outputPort_1_Daemon_CP_814_elements(111)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_814_elements(115);
      outputPort_1_Daemon_CP_814_elements(102) <= phi_mux_reqs(1);
      phi_stmt_608_phi_seq_1063 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_608_phi_seq_1063") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_814_elements(97), 
          phi_sample_ack => outputPort_1_Daemon_CP_814_elements(98), 
          phi_update_req => outputPort_1_Daemon_CP_814_elements(99), 
          phi_update_ack => outputPort_1_Daemon_CP_814_elements(100), 
          phi_mux_ack => outputPort_1_Daemon_CP_814_elements(105), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_613_phi_seq_1107_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_814_elements(124);
      outputPort_1_Daemon_CP_814_elements(127)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_814_elements(127);
      outputPort_1_Daemon_CP_814_elements(128)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_814_elements(129);
      outputPort_1_Daemon_CP_814_elements(125) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_814_elements(122);
      outputPort_1_Daemon_CP_814_elements(131)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_814_elements(133);
      outputPort_1_Daemon_CP_814_elements(132)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_814_elements(134);
      outputPort_1_Daemon_CP_814_elements(123) <= phi_mux_reqs(1);
      phi_stmt_613_phi_seq_1107 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_613_phi_seq_1107") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_814_elements(118), 
          phi_sample_ack => outputPort_1_Daemon_CP_814_elements(119), 
          phi_update_req => outputPort_1_Daemon_CP_814_elements(120), 
          phi_update_ack => outputPort_1_Daemon_CP_814_elements(121), 
          phi_mux_ack => outputPort_1_Daemon_CP_814_elements(126), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_617_phi_seq_1151_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_814_elements(143);
      outputPort_1_Daemon_CP_814_elements(146)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_814_elements(146);
      outputPort_1_Daemon_CP_814_elements(147)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_814_elements(148);
      outputPort_1_Daemon_CP_814_elements(144) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_814_elements(141);
      outputPort_1_Daemon_CP_814_elements(150)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_814_elements(152);
      outputPort_1_Daemon_CP_814_elements(151)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_814_elements(153);
      outputPort_1_Daemon_CP_814_elements(142) <= phi_mux_reqs(1);
      phi_stmt_617_phi_seq_1151 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_617_phi_seq_1151") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_814_elements(137), 
          phi_sample_ack => outputPort_1_Daemon_CP_814_elements(138), 
          phi_update_req => outputPort_1_Daemon_CP_814_elements(139), 
          phi_update_ack => outputPort_1_Daemon_CP_814_elements(140), 
          phi_mux_ack => outputPort_1_Daemon_CP_814_elements(145), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_839_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= outputPort_1_Daemon_CP_814_elements(7);
        preds(1)  <= outputPort_1_Daemon_CP_814_elements(8);
        entry_tmerge_839 : transition_merge -- 
          generic map(name => " entry_tmerge_839")
          port map (preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u3_u1_645_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_651_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_658_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_664_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_706_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_714_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_722_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_730_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_747_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_754_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_762_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_769_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_780_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_786_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_793_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_799_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_687_wire : std_logic_vector(0 downto 0);
    signal MUX_648_wire : std_logic_vector(0 downto 0);
    signal MUX_654_wire : std_logic_vector(0 downto 0);
    signal MUX_661_wire : std_logic_vector(0 downto 0);
    signal MUX_667_wire : std_logic_vector(0 downto 0);
    signal MUX_698_wire : std_logic_vector(7 downto 0);
    signal MUX_751_wire : std_logic_vector(31 downto 0);
    signal MUX_758_wire : std_logic_vector(31 downto 0);
    signal MUX_766_wire : std_logic_vector(31 downto 0);
    signal MUX_773_wire : std_logic_vector(31 downto 0);
    signal MUX_783_wire : std_logic_vector(0 downto 0);
    signal MUX_789_wire : std_logic_vector(0 downto 0);
    signal MUX_796_wire : std_logic_vector(0 downto 0);
    signal MUX_802_wire : std_logic_vector(0 downto 0);
    signal NEQ_u3_u1_684_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_703_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_711_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_719_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_727_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_655_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_668_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_790_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_803_wire : std_logic_vector(0 downto 0);
    signal OR_u32_u32_759_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_774_wire : std_logic_vector(31 downto 0);
    signal RPIPE_noblock_obuf_1_1_597_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_2_1_602_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_3_1_607_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_4_1_612_wire : std_logic_vector(32 downto 0);
    signal R_ONE_3_619_wire_constant : std_logic_vector(2 downto 0);
    signal R_ZERO_33_595_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_600_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_605_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_610_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_3_615_wire_constant : std_logic_vector(2 downto 0);
    signal R_ZERO_8_591_wire_constant : std_logic_vector(7 downto 0);
    signal SUB_u8_u8_696_wire : std_logic_vector(7 downto 0);
    signal active_packet_613 : std_logic_vector(2 downto 0);
    signal data_to_out_776 : std_logic_vector(31 downto 0);
    signal down_counter_589 : std_logic_vector(7 downto 0);
    signal konst_624_wire_constant : std_logic_vector(32 downto 0);
    signal konst_629_wire_constant : std_logic_vector(32 downto 0);
    signal konst_634_wire_constant : std_logic_vector(32 downto 0);
    signal konst_639_wire_constant : std_logic_vector(32 downto 0);
    signal konst_644_wire_constant : std_logic_vector(2 downto 0);
    signal konst_647_wire_constant : std_logic_vector(0 downto 0);
    signal konst_650_wire_constant : std_logic_vector(2 downto 0);
    signal konst_653_wire_constant : std_logic_vector(0 downto 0);
    signal konst_657_wire_constant : std_logic_vector(2 downto 0);
    signal konst_660_wire_constant : std_logic_vector(0 downto 0);
    signal konst_663_wire_constant : std_logic_vector(2 downto 0);
    signal konst_666_wire_constant : std_logic_vector(0 downto 0);
    signal konst_683_wire_constant : std_logic_vector(2 downto 0);
    signal konst_686_wire_constant : std_logic_vector(7 downto 0);
    signal konst_692_wire_constant : std_logic_vector(7 downto 0);
    signal konst_695_wire_constant : std_logic_vector(7 downto 0);
    signal konst_705_wire_constant : std_logic_vector(2 downto 0);
    signal konst_713_wire_constant : std_logic_vector(2 downto 0);
    signal konst_721_wire_constant : std_logic_vector(2 downto 0);
    signal konst_729_wire_constant : std_logic_vector(2 downto 0);
    signal konst_746_wire_constant : std_logic_vector(2 downto 0);
    signal konst_750_wire_constant : std_logic_vector(31 downto 0);
    signal konst_753_wire_constant : std_logic_vector(2 downto 0);
    signal konst_757_wire_constant : std_logic_vector(31 downto 0);
    signal konst_761_wire_constant : std_logic_vector(2 downto 0);
    signal konst_765_wire_constant : std_logic_vector(31 downto 0);
    signal konst_768_wire_constant : std_logic_vector(2 downto 0);
    signal konst_772_wire_constant : std_logic_vector(31 downto 0);
    signal konst_779_wire_constant : std_logic_vector(2 downto 0);
    signal konst_782_wire_constant : std_logic_vector(0 downto 0);
    signal konst_785_wire_constant : std_logic_vector(2 downto 0);
    signal konst_788_wire_constant : std_logic_vector(0 downto 0);
    signal konst_792_wire_constant : std_logic_vector(2 downto 0);
    signal konst_795_wire_constant : std_logic_vector(0 downto 0);
    signal konst_798_wire_constant : std_logic_vector(2 downto 0);
    signal konst_801_wire_constant : std_logic_vector(0 downto 0);
    signal konst_811_wire_constant : std_logic_vector(0 downto 0);
    signal next_active_packet_680 : std_logic_vector(2 downto 0);
    signal next_active_packet_680_616_buffered : std_logic_vector(2 downto 0);
    signal next_down_counter_700 : std_logic_vector(7 downto 0);
    signal next_down_counter_700_592_buffered : std_logic_vector(7 downto 0);
    signal next_pkt_priority_680 : std_logic_vector(2 downto 0);
    signal next_pkt_priority_680_620_buffered : std_logic_vector(2 downto 0);
    signal p1_valid_626 : std_logic_vector(0 downto 0);
    signal p2_valid_631 : std_logic_vector(0 downto 0);
    signal p3_valid_636 : std_logic_vector(0 downto 0);
    signal p4_valid_641 : std_logic_vector(0 downto 0);
    signal pkt_1_e_word_593 : std_logic_vector(32 downto 0);
    signal pkt_2_e_word_598 : std_logic_vector(32 downto 0);
    signal pkt_3_e_word_603 : std_logic_vector(32 downto 0);
    signal pkt_4_e_word_608 : std_logic_vector(32 downto 0);
    signal pkt_priority_617 : std_logic_vector(2 downto 0);
    signal read_from_1_708 : std_logic_vector(0 downto 0);
    signal read_from_2_716 : std_logic_vector(0 downto 0);
    signal read_from_3_724 : std_logic_vector(0 downto 0);
    signal read_from_4_732 : std_logic_vector(0 downto 0);
    signal send_flag_805 : std_logic_vector(0 downto 0);
    signal slice_749_wire : std_logic_vector(31 downto 0);
    signal slice_756_wire : std_logic_vector(31 downto 0);
    signal slice_764_wire : std_logic_vector(31 downto 0);
    signal slice_771_wire : std_logic_vector(31 downto 0);
    signal started_new_packet_689 : std_logic_vector(0 downto 0);
    signal valid_active_pkt_word_read_670 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_ONE_3_619_wire_constant <= "001";
    R_ZERO_33_595_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_600_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_605_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_610_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_3_615_wire_constant <= "000";
    R_ZERO_8_591_wire_constant <= "00000000";
    konst_624_wire_constant <= "000000000000000000000000000100000";
    konst_629_wire_constant <= "000000000000000000000000000100000";
    konst_634_wire_constant <= "000000000000000000000000000100000";
    konst_639_wire_constant <= "000000000000000000000000000100000";
    konst_644_wire_constant <= "001";
    konst_647_wire_constant <= "0";
    konst_650_wire_constant <= "010";
    konst_653_wire_constant <= "0";
    konst_657_wire_constant <= "011";
    konst_660_wire_constant <= "0";
    konst_663_wire_constant <= "100";
    konst_666_wire_constant <= "0";
    konst_683_wire_constant <= "000";
    konst_686_wire_constant <= "00000000";
    konst_692_wire_constant <= "00111111";
    konst_695_wire_constant <= "00000001";
    konst_705_wire_constant <= "001";
    konst_713_wire_constant <= "010";
    konst_721_wire_constant <= "011";
    konst_729_wire_constant <= "100";
    konst_746_wire_constant <= "001";
    konst_750_wire_constant <= "00000000000000000000000000000000";
    konst_753_wire_constant <= "010";
    konst_757_wire_constant <= "00000000000000000000000000000000";
    konst_761_wire_constant <= "011";
    konst_765_wire_constant <= "00000000000000000000000000000000";
    konst_768_wire_constant <= "100";
    konst_772_wire_constant <= "00000000000000000000000000000000";
    konst_779_wire_constant <= "001";
    konst_782_wire_constant <= "0";
    konst_785_wire_constant <= "010";
    konst_788_wire_constant <= "0";
    konst_792_wire_constant <= "011";
    konst_795_wire_constant <= "0";
    konst_798_wire_constant <= "100";
    konst_801_wire_constant <= "0";
    konst_811_wire_constant <= "1";
    phi_stmt_589: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_8_591_wire_constant & next_down_counter_700_592_buffered;
      req <= phi_stmt_589_req_0 & phi_stmt_589_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_589",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_589_ack_0,
          idata => idata,
          odata => down_counter_589,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_589
    phi_stmt_593: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_595_wire_constant & RPIPE_noblock_obuf_1_1_597_wire;
      req <= phi_stmt_593_req_0 & phi_stmt_593_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_593",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_593_ack_0,
          idata => idata,
          odata => pkt_1_e_word_593,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_593
    phi_stmt_598: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_600_wire_constant & RPIPE_noblock_obuf_2_1_602_wire;
      req <= phi_stmt_598_req_0 & phi_stmt_598_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_598",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_598_ack_0,
          idata => idata,
          odata => pkt_2_e_word_598,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_598
    phi_stmt_603: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_605_wire_constant & RPIPE_noblock_obuf_3_1_607_wire;
      req <= phi_stmt_603_req_0 & phi_stmt_603_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_603",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_603_ack_0,
          idata => idata,
          odata => pkt_3_e_word_603,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_603
    phi_stmt_608: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_610_wire_constant & RPIPE_noblock_obuf_4_1_612_wire;
      req <= phi_stmt_608_req_0 & phi_stmt_608_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_608",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_608_ack_0,
          idata => idata,
          odata => pkt_4_e_word_608,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_608
    phi_stmt_613: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_3_615_wire_constant & next_active_packet_680_616_buffered;
      req <= phi_stmt_613_req_0 & phi_stmt_613_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_613",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_613_ack_0,
          idata => idata,
          odata => active_packet_613,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_613
    phi_stmt_617: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ONE_3_619_wire_constant & next_pkt_priority_680_620_buffered;
      req <= phi_stmt_617_req_0 & phi_stmt_617_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_617",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_617_ack_0,
          idata => idata,
          odata => pkt_priority_617,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_617
    -- flow-through select operator MUX_648_inst
    MUX_648_wire <= p1_valid_626 when (EQ_u3_u1_645_wire(0) /=  '0') else konst_647_wire_constant;
    -- flow-through select operator MUX_654_inst
    MUX_654_wire <= p2_valid_631 when (EQ_u3_u1_651_wire(0) /=  '0') else konst_653_wire_constant;
    -- flow-through select operator MUX_661_inst
    MUX_661_wire <= p3_valid_636 when (EQ_u3_u1_658_wire(0) /=  '0') else konst_660_wire_constant;
    -- flow-through select operator MUX_667_inst
    MUX_667_wire <= p4_valid_641 when (EQ_u3_u1_664_wire(0) /=  '0') else konst_666_wire_constant;
    -- flow-through select operator MUX_698_inst
    MUX_698_wire <= SUB_u8_u8_696_wire when (valid_active_pkt_word_read_670(0) /=  '0') else down_counter_589;
    -- flow-through select operator MUX_699_inst
    next_down_counter_700 <= konst_692_wire_constant when (started_new_packet_689(0) /=  '0') else MUX_698_wire;
    -- flow-through select operator MUX_751_inst
    MUX_751_wire <= slice_749_wire when (EQ_u3_u1_747_wire(0) /=  '0') else konst_750_wire_constant;
    -- flow-through select operator MUX_758_inst
    MUX_758_wire <= slice_756_wire when (EQ_u3_u1_754_wire(0) /=  '0') else konst_757_wire_constant;
    -- flow-through select operator MUX_766_inst
    MUX_766_wire <= slice_764_wire when (EQ_u3_u1_762_wire(0) /=  '0') else konst_765_wire_constant;
    -- flow-through select operator MUX_773_inst
    MUX_773_wire <= slice_771_wire when (EQ_u3_u1_769_wire(0) /=  '0') else konst_772_wire_constant;
    -- flow-through select operator MUX_783_inst
    MUX_783_wire <= p1_valid_626 when (EQ_u3_u1_780_wire(0) /=  '0') else konst_782_wire_constant;
    -- flow-through select operator MUX_789_inst
    MUX_789_wire <= p2_valid_631 when (EQ_u3_u1_786_wire(0) /=  '0') else konst_788_wire_constant;
    -- flow-through select operator MUX_796_inst
    MUX_796_wire <= p3_valid_636 when (EQ_u3_u1_793_wire(0) /=  '0') else konst_795_wire_constant;
    -- flow-through select operator MUX_802_inst
    MUX_802_wire <= p4_valid_641 when (EQ_u3_u1_799_wire(0) /=  '0') else konst_801_wire_constant;
    -- flow-through slice operator slice_749_inst
    slice_749_wire <= pkt_1_e_word_593(31 downto 0);
    -- flow-through slice operator slice_756_inst
    slice_756_wire <= pkt_2_e_word_598(31 downto 0);
    -- flow-through slice operator slice_764_inst
    slice_764_wire <= pkt_3_e_word_603(31 downto 0);
    -- flow-through slice operator slice_771_inst
    slice_771_wire <= pkt_4_e_word_608(31 downto 0);
    next_active_packet_680_616_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_active_packet_680_616_buf_req_0;
      next_active_packet_680_616_buf_ack_0<= wack(0);
      rreq(0) <= next_active_packet_680_616_buf_req_1;
      next_active_packet_680_616_buf_ack_1<= rack(0);
      next_active_packet_680_616_buf : InterlockBuffer generic map ( -- 
        name => "next_active_packet_680_616_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_active_packet_680,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_active_packet_680_616_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_down_counter_700_592_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_down_counter_700_592_buf_req_0;
      next_down_counter_700_592_buf_ack_0<= wack(0);
      rreq(0) <= next_down_counter_700_592_buf_req_1;
      next_down_counter_700_592_buf_ack_1<= rack(0);
      next_down_counter_700_592_buf : InterlockBuffer generic map ( -- 
        name => "next_down_counter_700_592_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_down_counter_700,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_down_counter_700_592_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_pkt_priority_680_620_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_pkt_priority_680_620_buf_req_0;
      next_pkt_priority_680_620_buf_ack_0<= wack(0);
      rreq(0) <= next_pkt_priority_680_620_buf_req_1;
      next_pkt_priority_680_620_buf_ack_1<= rack(0);
      next_pkt_priority_680_620_buf : InterlockBuffer generic map ( -- 
        name => "next_pkt_priority_680_620_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_pkt_priority_680,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_pkt_priority_680_620_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_587_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_811_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_587_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_587_branch_req_0,
          ack0 => do_while_stmt_587_branch_ack_0,
          ack1 => do_while_stmt_587_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator AND_u1_u1_688_inst
    process(NEQ_u3_u1_684_wire, EQ_u8_u1_687_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NEQ_u3_u1_684_wire, EQ_u8_u1_687_wire, tmp_var);
      started_new_packet_689 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_625_inst
    process(pkt_1_e_word_593) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_1_e_word_593, konst_624_wire_constant, tmp_var);
      p1_valid_626 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_630_inst
    process(pkt_2_e_word_598) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_2_e_word_598, konst_629_wire_constant, tmp_var);
      p2_valid_631 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_635_inst
    process(pkt_3_e_word_603) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_3_e_word_603, konst_634_wire_constant, tmp_var);
      p3_valid_636 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_640_inst
    process(pkt_4_e_word_608) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_4_e_word_608, konst_639_wire_constant, tmp_var);
      p4_valid_641 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_645_inst
    process(active_packet_613) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_613, konst_644_wire_constant, tmp_var);
      EQ_u3_u1_645_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_651_inst
    process(active_packet_613) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_613, konst_650_wire_constant, tmp_var);
      EQ_u3_u1_651_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_658_inst
    process(active_packet_613) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_613, konst_657_wire_constant, tmp_var);
      EQ_u3_u1_658_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_664_inst
    process(active_packet_613) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_613, konst_663_wire_constant, tmp_var);
      EQ_u3_u1_664_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_706_inst
    process(next_active_packet_680) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_680, konst_705_wire_constant, tmp_var);
      EQ_u3_u1_706_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_714_inst
    process(next_active_packet_680) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_680, konst_713_wire_constant, tmp_var);
      EQ_u3_u1_714_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_722_inst
    process(next_active_packet_680) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_680, konst_721_wire_constant, tmp_var);
      EQ_u3_u1_722_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_730_inst
    process(next_active_packet_680) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_680, konst_729_wire_constant, tmp_var);
      EQ_u3_u1_730_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_747_inst
    process(next_active_packet_680) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_680, konst_746_wire_constant, tmp_var);
      EQ_u3_u1_747_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_754_inst
    process(next_active_packet_680) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_680, konst_753_wire_constant, tmp_var);
      EQ_u3_u1_754_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_762_inst
    process(next_active_packet_680) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_680, konst_761_wire_constant, tmp_var);
      EQ_u3_u1_762_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_769_inst
    process(next_active_packet_680) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_680, konst_768_wire_constant, tmp_var);
      EQ_u3_u1_769_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_780_inst
    process(next_active_packet_680) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_680, konst_779_wire_constant, tmp_var);
      EQ_u3_u1_780_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_786_inst
    process(next_active_packet_680) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_680, konst_785_wire_constant, tmp_var);
      EQ_u3_u1_786_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_793_inst
    process(next_active_packet_680) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_680, konst_792_wire_constant, tmp_var);
      EQ_u3_u1_793_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_799_inst
    process(next_active_packet_680) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_680, konst_798_wire_constant, tmp_var);
      EQ_u3_u1_799_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_687_inst
    process(down_counter_589) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(down_counter_589, konst_686_wire_constant, tmp_var);
      EQ_u8_u1_687_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u3_u1_684_inst
    process(next_active_packet_680) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(next_active_packet_680, konst_683_wire_constant, tmp_var);
      NEQ_u3_u1_684_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_703_inst
    process(p1_valid_626) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_626, tmp_var);
      NOT_u1_u1_703_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_711_inst
    process(p2_valid_631) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_631, tmp_var);
      NOT_u1_u1_711_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_719_inst
    process(p3_valid_636) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_636, tmp_var);
      NOT_u1_u1_719_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_727_inst
    process(p4_valid_641) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_641, tmp_var);
      NOT_u1_u1_727_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_655_inst
    process(MUX_648_wire, MUX_654_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_648_wire, MUX_654_wire, tmp_var);
      OR_u1_u1_655_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_668_inst
    process(MUX_661_wire, MUX_667_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_661_wire, MUX_667_wire, tmp_var);
      OR_u1_u1_668_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_669_inst
    process(OR_u1_u1_655_wire, OR_u1_u1_668_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_655_wire, OR_u1_u1_668_wire, tmp_var);
      valid_active_pkt_word_read_670 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_707_inst
    process(NOT_u1_u1_703_wire, EQ_u3_u1_706_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_703_wire, EQ_u3_u1_706_wire, tmp_var);
      read_from_1_708 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_715_inst
    process(NOT_u1_u1_711_wire, EQ_u3_u1_714_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_711_wire, EQ_u3_u1_714_wire, tmp_var);
      read_from_2_716 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_723_inst
    process(NOT_u1_u1_719_wire, EQ_u3_u1_722_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_719_wire, EQ_u3_u1_722_wire, tmp_var);
      read_from_3_724 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_731_inst
    process(NOT_u1_u1_727_wire, EQ_u3_u1_730_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_727_wire, EQ_u3_u1_730_wire, tmp_var);
      read_from_4_732 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_790_inst
    process(MUX_783_wire, MUX_789_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_783_wire, MUX_789_wire, tmp_var);
      OR_u1_u1_790_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_803_inst
    process(MUX_796_wire, MUX_802_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_796_wire, MUX_802_wire, tmp_var);
      OR_u1_u1_803_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_804_inst
    process(OR_u1_u1_790_wire, OR_u1_u1_803_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_790_wire, OR_u1_u1_803_wire, tmp_var);
      send_flag_805 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_759_inst
    process(MUX_751_wire, MUX_758_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_751_wire, MUX_758_wire, tmp_var);
      OR_u32_u32_759_wire <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_774_inst
    process(MUX_766_wire, MUX_773_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_766_wire, MUX_773_wire, tmp_var);
      OR_u32_u32_774_wire <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_775_inst
    process(OR_u32_u32_759_wire, OR_u32_u32_774_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u32_u32_759_wire, OR_u32_u32_774_wire, tmp_var);
      data_to_out_776 <= tmp_var; --
    end process;
    -- binary operator SUB_u8_u8_696_inst
    process(down_counter_589) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSub_proc(down_counter_589, konst_695_wire_constant, tmp_var);
      SUB_u8_u8_696_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_noblock_obuf_1_1_597_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_1_1_597_inst_req_0;
      RPIPE_noblock_obuf_1_1_597_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_1_1_597_inst_req_1;
      RPIPE_noblock_obuf_1_1_597_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_1_708(0);
      RPIPE_noblock_obuf_1_1_597_wire <= data_out(32 downto 0);
      noblock_obuf_1_1_read_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_1_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_1_read_0: InputPortRevised -- 
        generic map ( name => "noblock_obuf_1_1_read_0", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_1_1_pipe_read_req(0),
          oack => noblock_obuf_1_1_pipe_read_ack(0),
          odata => noblock_obuf_1_1_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_noblock_obuf_2_1_602_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_2_1_602_inst_req_0;
      RPIPE_noblock_obuf_2_1_602_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_2_1_602_inst_req_1;
      RPIPE_noblock_obuf_2_1_602_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_2_716(0);
      RPIPE_noblock_obuf_2_1_602_wire <= data_out(32 downto 0);
      noblock_obuf_2_1_read_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_1_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_1_read_1: InputPortRevised -- 
        generic map ( name => "noblock_obuf_2_1_read_1", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_2_1_pipe_read_req(0),
          oack => noblock_obuf_2_1_pipe_read_ack(0),
          odata => noblock_obuf_2_1_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_noblock_obuf_3_1_607_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_3_1_607_inst_req_0;
      RPIPE_noblock_obuf_3_1_607_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_3_1_607_inst_req_1;
      RPIPE_noblock_obuf_3_1_607_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_3_724(0);
      RPIPE_noblock_obuf_3_1_607_wire <= data_out(32 downto 0);
      noblock_obuf_3_1_read_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_1_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_1_read_2: InputPortRevised -- 
        generic map ( name => "noblock_obuf_3_1_read_2", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_3_1_pipe_read_req(0),
          oack => noblock_obuf_3_1_pipe_read_ack(0),
          odata => noblock_obuf_3_1_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_noblock_obuf_4_1_612_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_4_1_612_inst_req_0;
      RPIPE_noblock_obuf_4_1_612_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_4_1_612_inst_req_1;
      RPIPE_noblock_obuf_4_1_612_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_4_732(0);
      RPIPE_noblock_obuf_4_1_612_wire <= data_out(32 downto 0);
      noblock_obuf_4_1_read_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_1_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_1_read_3: InputPortRevised -- 
        generic map ( name => "noblock_obuf_4_1_read_3", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_4_1_pipe_read_req(0),
          oack => noblock_obuf_4_1_pipe_read_ack(0),
          odata => noblock_obuf_4_1_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_out_data_1_807_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_out_data_1_807_inst_req_0;
      WPIPE_out_data_1_807_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_out_data_1_807_inst_req_1;
      WPIPE_out_data_1_807_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_flag_805(0);
      data_in <= data_to_out_776;
      out_data_1_write_0_gI: SplitGuardInterface generic map(name => "out_data_1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      out_data_1_write_0: OutputPortRevised -- 
        generic map ( name => "out_data_1", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => out_data_1_pipe_write_req(0),
          oack => out_data_1_pipe_write_ack(0),
          odata => out_data_1_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    volatile_operator_prioritySelect_1874: prioritySelect_Volatile port map(down_counter => down_counter_589, active_packet => active_packet_613, pkt_priority => pkt_priority_617, p1_valid => p1_valid_626, p2_valid => p2_valid_631, p3_valid => p3_valid_636, p4_valid => p4_valid_641, next_active_packet => next_active_packet_680, next_pkt_priority => next_pkt_priority_680); 
    -- 
  end Block; -- data_path
  -- 
end outputPort_1_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity outputPort_2_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    noblock_obuf_1_2_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_2_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_3_2_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_2_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_4_2_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_2_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_2_2_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_2_pipe_read_data : in   std_logic_vector(32 downto 0);
    out_data_2_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_2_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity outputPort_2_Daemon;
architecture outputPort_2_Daemon_arch of outputPort_2_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal outputPort_2_Daemon_CP_1176_start: Boolean;
  signal outputPort_2_Daemon_CP_1176_symbol: Boolean;
  -- volatile/operator module components. 
  component prioritySelect_Volatile is -- 
    port ( -- 
      down_counter : in  std_logic_vector(7 downto 0);
      active_packet : in  std_logic_vector(2 downto 0);
      pkt_priority : in  std_logic_vector(2 downto 0);
      p1_valid : in  std_logic_vector(0 downto 0);
      p2_valid : in  std_logic_vector(0 downto 0);
      p3_valid : in  std_logic_vector(0 downto 0);
      p4_valid : in  std_logic_vector(0 downto 0);
      next_active_packet : out  std_logic_vector(2 downto 0);
      next_pkt_priority : out  std_logic_vector(2 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal do_while_stmt_816_branch_ack_1 : boolean;
  signal next_active_packet_909_845_buf_req_1 : boolean;
  signal next_active_packet_909_845_buf_req_0 : boolean;
  signal WPIPE_out_data_2_1036_inst_ack_0 : boolean;
  signal next_active_packet_909_845_buf_ack_0 : boolean;
  signal next_pkt_priority_909_849_buf_req_0 : boolean;
  signal next_pkt_priority_909_849_buf_ack_0 : boolean;
  signal next_active_packet_909_845_buf_ack_1 : boolean;
  signal next_pkt_priority_909_849_buf_ack_1 : boolean;
  signal phi_stmt_842_req_0 : boolean;
  signal next_pkt_priority_909_849_buf_req_1 : boolean;
  signal phi_stmt_842_req_1 : boolean;
  signal phi_stmt_846_req_0 : boolean;
  signal phi_stmt_818_req_1 : boolean;
  signal do_while_stmt_816_branch_req_0 : boolean;
  signal phi_stmt_818_req_0 : boolean;
  signal phi_stmt_846_ack_0 : boolean;
  signal phi_stmt_846_req_1 : boolean;
  signal WPIPE_out_data_2_1036_inst_req_1 : boolean;
  signal phi_stmt_842_ack_0 : boolean;
  signal WPIPE_out_data_2_1036_inst_ack_1 : boolean;
  signal do_while_stmt_816_branch_ack_0 : boolean;
  signal WPIPE_out_data_2_1036_inst_req_0 : boolean;
  signal phi_stmt_818_ack_0 : boolean;
  signal next_down_counter_929_821_buf_req_0 : boolean;
  signal next_down_counter_929_821_buf_ack_0 : boolean;
  signal next_down_counter_929_821_buf_req_1 : boolean;
  signal next_down_counter_929_821_buf_ack_1 : boolean;
  signal phi_stmt_822_req_1 : boolean;
  signal phi_stmt_822_req_0 : boolean;
  signal phi_stmt_822_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_2_826_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_1_2_826_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_2_826_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_1_2_826_inst_ack_1 : boolean;
  signal phi_stmt_827_req_1 : boolean;
  signal phi_stmt_827_req_0 : boolean;
  signal phi_stmt_827_ack_0 : boolean;
  signal RPIPE_noblock_obuf_2_2_831_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_2_2_831_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_2_2_831_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_2_2_831_inst_ack_1 : boolean;
  signal phi_stmt_832_req_1 : boolean;
  signal phi_stmt_832_req_0 : boolean;
  signal phi_stmt_832_ack_0 : boolean;
  signal RPIPE_noblock_obuf_3_2_836_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_3_2_836_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_3_2_836_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_3_2_836_inst_ack_1 : boolean;
  signal phi_stmt_837_req_1 : boolean;
  signal phi_stmt_837_req_0 : boolean;
  signal phi_stmt_837_ack_0 : boolean;
  signal RPIPE_noblock_obuf_4_2_841_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_4_2_841_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_4_2_841_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_4_2_841_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "outputPort_2_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  outputPort_2_Daemon_CP_1176_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "outputPort_2_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_2_Daemon_CP_1176_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= outputPort_2_Daemon_CP_1176_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_2_Daemon_CP_1176_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  outputPort_2_Daemon_CP_1176: Block -- control-path 
    signal outputPort_2_Daemon_CP_1176_elements: BooleanArray(161 downto 0);
    -- 
  begin -- 
    outputPort_2_Daemon_CP_1176_elements(0) <= outputPort_2_Daemon_CP_1176_start;
    outputPort_2_Daemon_CP_1176_symbol <= outputPort_2_Daemon_CP_1176_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_815/branch_block_stmt_815__entry__
      -- CP-element group 0: 	 branch_block_stmt_815/$entry
      -- CP-element group 0: 	 branch_block_stmt_815/do_while_stmt_816__entry__
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	161 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_815/branch_block_stmt_815__exit__
      -- CP-element group 1: 	 branch_block_stmt_815/$exit
      -- CP-element group 1: 	 branch_block_stmt_815/do_while_stmt_816__exit__
      -- 
    outputPort_2_Daemon_CP_1176_elements(1) <= outputPort_2_Daemon_CP_1176_elements(161);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816__entry__
      -- CP-element group 2: 	 branch_block_stmt_815/do_while_stmt_816/$entry
      -- 
    outputPort_2_Daemon_CP_1176_elements(2) <= outputPort_2_Daemon_CP_1176_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	161 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816__exit__
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_815/do_while_stmt_816/loop_back
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	159 
    -- CP-element group 5: 	160 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_815/do_while_stmt_816/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_815/do_while_stmt_816/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_815/do_while_stmt_816/condition_done
      -- 
    outputPort_2_Daemon_CP_1176_elements(5) <= outputPort_2_Daemon_CP_1176_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	158 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_815/do_while_stmt_816/loop_body_done
      -- 
    outputPort_2_Daemon_CP_1176_elements(6) <= outputPort_2_Daemon_CP_1176_elements(158);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	141 
    -- CP-element group 7: 	21 
    -- CP-element group 7: 	40 
    -- CP-element group 7: 	61 
    -- CP-element group 7: 	82 
    -- CP-element group 7: 	103 
    -- CP-element group 7: 	124 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/back_edge_to_loop_body
      -- 
    outputPort_2_Daemon_CP_1176_elements(7) <= outputPort_2_Daemon_CP_1176_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	143 
    -- CP-element group 8: 	23 
    -- CP-element group 8: 	42 
    -- CP-element group 8: 	63 
    -- CP-element group 8: 	84 
    -- CP-element group 8: 	105 
    -- CP-element group 8: 	126 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/first_time_through_loop_body
      -- 
    outputPort_2_Daemon_CP_1176_elements(8) <= outputPort_2_Daemon_CP_1176_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	157 
    -- CP-element group 9: 	138 
    -- CP-element group 9: 	137 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	34 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	55 
    -- CP-element group 9: 	56 
    -- CP-element group 9: 	76 
    -- CP-element group 9: 	77 
    -- CP-element group 9: 	97 
    -- CP-element group 9: 	98 
    -- CP-element group 9: 	118 
    -- CP-element group 9: 	119 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/$entry
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	157 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/condition_evaluated
      -- 
    condition_evaluated_1200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(10), ack => do_while_stmt_816_branch_req_0); -- 
    outputPort_2_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(157) & outputPort_2_Daemon_CP_1176_elements(14);
      gj_outputPort_2_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	137 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	55 
    -- CP-element group 11: 	76 
    -- CP-element group 11: 	97 
    -- CP-element group 11: 	118 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	57 
    -- CP-element group 11: 	78 
    -- CP-element group 11: 	99 
    -- CP-element group 11: 	120 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_846_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/aggregated_phi_sample_req
      -- 
    outputPort_2_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(137) & outputPort_2_Daemon_CP_1176_elements(15) & outputPort_2_Daemon_CP_1176_elements(34) & outputPort_2_Daemon_CP_1176_elements(55) & outputPort_2_Daemon_CP_1176_elements(76) & outputPort_2_Daemon_CP_1176_elements(97) & outputPort_2_Daemon_CP_1176_elements(118) & outputPort_2_Daemon_CP_1176_elements(14);
      gj_outputPort_2_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	139 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	37 
    -- CP-element group 12: 	58 
    -- CP-element group 12: 	79 
    -- CP-element group 12: 	100 
    -- CP-element group 12: 	121 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	158 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	137 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	34 
    -- CP-element group 12: 	55 
    -- CP-element group 12: 	76 
    -- CP-element group 12: 	97 
    -- CP-element group 12: 	118 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_846_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_818_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_842_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_822_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_827_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_832_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_837_sample_completed_
      -- 
    outputPort_2_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(139) & outputPort_2_Daemon_CP_1176_elements(18) & outputPort_2_Daemon_CP_1176_elements(37) & outputPort_2_Daemon_CP_1176_elements(58) & outputPort_2_Daemon_CP_1176_elements(79) & outputPort_2_Daemon_CP_1176_elements(100) & outputPort_2_Daemon_CP_1176_elements(121);
      gj_outputPort_2_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	138 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	35 
    -- CP-element group 13: 	56 
    -- CP-element group 13: 	77 
    -- CP-element group 13: 	98 
    -- CP-element group 13: 	119 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	19 
    -- CP-element group 13: 	38 
    -- CP-element group 13: 	59 
    -- CP-element group 13: 	80 
    -- CP-element group 13: 	101 
    -- CP-element group 13: 	122 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_846_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/aggregated_phi_update_req
      -- 
    outputPort_2_Daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(138) & outputPort_2_Daemon_CP_1176_elements(16) & outputPort_2_Daemon_CP_1176_elements(35) & outputPort_2_Daemon_CP_1176_elements(56) & outputPort_2_Daemon_CP_1176_elements(77) & outputPort_2_Daemon_CP_1176_elements(98) & outputPort_2_Daemon_CP_1176_elements(119);
      gj_outputPort_2_Daemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	140 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	60 
    -- CP-element group 14: 	81 
    -- CP-element group 14: 	102 
    -- CP-element group 14: 	123 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/aggregated_phi_update_ack
      -- 
    outputPort_2_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(140) & outputPort_2_Daemon_CP_1176_elements(20) & outputPort_2_Daemon_CP_1176_elements(39) & outputPort_2_Daemon_CP_1176_elements(60) & outputPort_2_Daemon_CP_1176_elements(81) & outputPort_2_Daemon_CP_1176_elements(102) & outputPort_2_Daemon_CP_1176_elements(123);
      gj_outputPort_2_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_818_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	155 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_818_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(155);
      gj_outputPort_2_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_818_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(17) <= outputPort_2_Daemon_CP_1176_elements(11);
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_818_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_818_update_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(19) <= outputPort_2_Daemon_CP_1176_elements(13);
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	154 
    -- CP-element group 20: 	14 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_818_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_818_update_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_818_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(21) <= outputPort_2_Daemon_CP_1176_elements(7);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_818_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_818_loopback_sample_req_ps
      -- 
    phi_stmt_818_loopback_sample_req_1215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_818_loopback_sample_req_1215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(22), ack => phi_stmt_818_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_818_entry_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(23) <= outputPort_2_Daemon_CP_1176_elements(8);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_818_entry_sample_req
      -- CP-element group 24: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_818_entry_sample_req_ps
      -- 
    phi_stmt_818_entry_sample_req_1218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_818_entry_sample_req_1218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(24), ack => phi_stmt_818_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_818_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_818_phi_mux_ack_ps
      -- 
    phi_stmt_818_phi_mux_ack_1221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_818_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_8_820_sample_start__ps
      -- CP-element group 26: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_8_820_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_8_820_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_8_820_sample_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_8_820_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_8_820_update_start_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_8_820_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(28) <= outputPort_2_Daemon_CP_1176_elements(29);
    -- CP-element group 29:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	28 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_8_820_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(29) is a control-delay.
    cp_element_29_delay: control_delay_element  generic map(name => " 29_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_1176_elements(27), ack => outputPort_2_Daemon_CP_1176_elements(29), clk => clk, reset =>reset);
    -- CP-element group 30:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_down_counter_821_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_down_counter_821_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_down_counter_821_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_down_counter_821_Sample/req
      -- 
    req_1242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(30), ack => next_down_counter_929_821_buf_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_down_counter_821_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_down_counter_821_update_start_
      -- CP-element group 31: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_down_counter_821_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_down_counter_821_Update/req
      -- 
    req_1247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(31), ack => next_down_counter_929_821_buf_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_down_counter_821_sample_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_down_counter_821_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_down_counter_821_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_down_counter_821_Sample/ack
      -- 
    ack_1243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_929_821_buf_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(32)); -- 
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_down_counter_821_update_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_down_counter_821_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_down_counter_821_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_down_counter_821_Update/ack
      -- 
    ack_1248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_929_821_buf_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(33)); -- 
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	9 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	12 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	11 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_822_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	155 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	13 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_822_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(155);
      gj_outputPort_2_Daemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	11 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_822_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(36) <= outputPort_2_Daemon_CP_1176_elements(11);
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	12 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_822_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_822_update_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(38) <= outputPort_2_Daemon_CP_1176_elements(13);
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	154 
    -- CP-element group 39: 	14 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_822_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_822_update_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	7 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_822_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(40) <= outputPort_2_Daemon_CP_1176_elements(7);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_822_loopback_sample_req
      -- CP-element group 41: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_822_loopback_sample_req_ps
      -- 
    phi_stmt_822_loopback_sample_req_1259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_822_loopback_sample_req_1259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(41), ack => phi_stmt_822_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	8 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_822_entry_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(42) <= outputPort_2_Daemon_CP_1176_elements(8);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_822_entry_sample_req
      -- CP-element group 43: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_822_entry_sample_req_ps
      -- 
    phi_stmt_822_entry_sample_req_1262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_822_entry_sample_req_1262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(43), ack => phi_stmt_822_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_822_phi_mux_ack
      -- CP-element group 44: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_822_phi_mux_ack_ps
      -- 
    phi_stmt_822_phi_mux_ack_1265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_822_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_824_sample_start__ps
      -- CP-element group 45: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_824_sample_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_824_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_824_sample_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_824_update_start__ps
      -- CP-element group 46: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_824_update_start_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_824_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(47) <= outputPort_2_Daemon_CP_1176_elements(48);
    -- CP-element group 48:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	47 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_824_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(48) is a control-delay.
    cp_element_48_delay: control_delay_element  generic map(name => " 48_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_1176_elements(46), ack => outputPort_2_Daemon_CP_1176_elements(48), clk => clk, reset =>reset);
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_1_2_826_sample_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_1_2_826_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	54 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_1_2_826_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_1_2_826_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_1_2_826_Sample/rr
      -- 
    rr_1286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(51), ack => RPIPE_noblock_obuf_1_2_826_inst_req_0); -- 
    outputPort_2_Daemon_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(49) & outputPort_2_Daemon_CP_1176_elements(54);
      gj_outputPort_2_Daemon_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: 	53 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_1_2_826_update_start_
      -- CP-element group 52: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_1_2_826_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_1_2_826_Update/cr
      -- 
    cr_1291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(52), ack => RPIPE_noblock_obuf_1_2_826_inst_req_1); -- 
    outputPort_2_Daemon_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(50) & outputPort_2_Daemon_CP_1176_elements(53);
      gj_outputPort_2_Daemon_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	52 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_1_2_826_sample_completed__ps
      -- CP-element group 53: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_1_2_826_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_1_2_826_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_1_2_826_Sample/ra
      -- 
    ra_1287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_2_826_inst_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(53)); -- 
    -- CP-element group 54:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	51 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_1_2_826_update_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_1_2_826_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_1_2_826_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_1_2_826_Update/ca
      -- 
    ca_1292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_2_826_inst_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(54)); -- 
    -- CP-element group 55:  join  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	9 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	12 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	11 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_827_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	9 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	155 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	13 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_827_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(155);
      gj_outputPort_2_Daemon_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	11 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_827_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(57) <= outputPort_2_Daemon_CP_1176_elements(11);
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	12 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_827_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	13 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_827_update_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(59) <= outputPort_2_Daemon_CP_1176_elements(13);
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	154 
    -- CP-element group 60: 	14 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_827_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_827_update_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	7 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_827_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(61) <= outputPort_2_Daemon_CP_1176_elements(7);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_827_loopback_sample_req
      -- CP-element group 62: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_827_loopback_sample_req_ps
      -- 
    phi_stmt_827_loopback_sample_req_1303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_827_loopback_sample_req_1303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(62), ack => phi_stmt_827_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	8 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_827_entry_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(63) <= outputPort_2_Daemon_CP_1176_elements(8);
    -- CP-element group 64:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_827_entry_sample_req
      -- CP-element group 64: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_827_entry_sample_req_ps
      -- 
    phi_stmt_827_entry_sample_req_1306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_827_entry_sample_req_1306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(64), ack => phi_stmt_827_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_827_phi_mux_ack
      -- CP-element group 65: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_827_phi_mux_ack_ps
      -- 
    phi_stmt_827_phi_mux_ack_1309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_827_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(65)); -- 
    -- CP-element group 66:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_829_sample_start__ps
      -- CP-element group 66: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_829_sample_completed__ps
      -- CP-element group 66: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_829_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_829_sample_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_829_update_start__ps
      -- CP-element group 67: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_829_update_start_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_829_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(68) <= outputPort_2_Daemon_CP_1176_elements(69);
    -- CP-element group 69:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	68 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_829_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(69) is a control-delay.
    cp_element_69_delay: control_delay_element  generic map(name => " 69_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_1176_elements(67), ack => outputPort_2_Daemon_CP_1176_elements(69), clk => clk, reset =>reset);
    -- CP-element group 70:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_2_2_831_sample_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(70) is bound as output of CP function.
    -- CP-element group 71:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_2_2_831_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: marked-predecessors 
    -- CP-element group 72: 	75 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_2_2_831_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_2_2_831_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_2_2_831_Sample/rr
      -- 
    rr_1330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(72), ack => RPIPE_noblock_obuf_2_2_831_inst_req_0); -- 
    outputPort_2_Daemon_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(70) & outputPort_2_Daemon_CP_1176_elements(75);
      gj_outputPort_2_Daemon_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: 	74 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_2_2_831_update_start_
      -- CP-element group 73: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_2_2_831_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_2_2_831_Update/cr
      -- 
    cr_1335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(73), ack => RPIPE_noblock_obuf_2_2_831_inst_req_1); -- 
    outputPort_2_Daemon_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(71) & outputPort_2_Daemon_CP_1176_elements(74);
      gj_outputPort_2_Daemon_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	73 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_2_2_831_sample_completed__ps
      -- CP-element group 74: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_2_2_831_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_2_2_831_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_2_2_831_Sample/ra
      -- 
    ra_1331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_2_831_inst_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(74)); -- 
    -- CP-element group 75:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	72 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_2_2_831_update_completed__ps
      -- CP-element group 75: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_2_2_831_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_2_2_831_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_2_2_831_Update/ca
      -- 
    ca_1336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_2_831_inst_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(75)); -- 
    -- CP-element group 76:  join  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	9 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	12 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	11 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_832_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	9 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	155 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	13 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_832_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(155);
      gj_outputPort_2_Daemon_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	11 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_832_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(78) <= outputPort_2_Daemon_CP_1176_elements(11);
    -- CP-element group 79:  join  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	12 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_832_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	13 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_832_update_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(80) <= outputPort_2_Daemon_CP_1176_elements(13);
    -- CP-element group 81:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	154 
    -- CP-element group 81: 	14 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_832_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_832_update_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	7 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_832_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(82) <= outputPort_2_Daemon_CP_1176_elements(7);
    -- CP-element group 83:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_832_loopback_sample_req
      -- CP-element group 83: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_832_loopback_sample_req_ps
      -- 
    phi_stmt_832_loopback_sample_req_1347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_832_loopback_sample_req_1347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(83), ack => phi_stmt_832_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(83) is bound as output of CP function.
    -- CP-element group 84:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	8 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_832_entry_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(84) <= outputPort_2_Daemon_CP_1176_elements(8);
    -- CP-element group 85:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_832_entry_sample_req
      -- CP-element group 85: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_832_entry_sample_req_ps
      -- 
    phi_stmt_832_entry_sample_req_1350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_832_entry_sample_req_1350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(85), ack => phi_stmt_832_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_832_phi_mux_ack_ps
      -- CP-element group 86: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_832_phi_mux_ack
      -- 
    phi_stmt_832_phi_mux_ack_1353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_832_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(86)); -- 
    -- CP-element group 87:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_834_sample_start__ps
      -- CP-element group 87: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_834_sample_completed__ps
      -- CP-element group 87: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_834_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_834_sample_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_834_update_start__ps
      -- CP-element group 88: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_834_update_start_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	90 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_834_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(89) <= outputPort_2_Daemon_CP_1176_elements(90);
    -- CP-element group 90:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	89 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_834_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(90) is a control-delay.
    cp_element_90_delay: control_delay_element  generic map(name => " 90_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_1176_elements(88), ack => outputPort_2_Daemon_CP_1176_elements(90), clk => clk, reset =>reset);
    -- CP-element group 91:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_3_2_836_sample_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(91) is bound as output of CP function.
    -- CP-element group 92:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_3_2_836_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(92) is bound as output of CP function.
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	96 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_3_2_836_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_3_2_836_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_3_2_836_Sample/rr
      -- 
    rr_1374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(93), ack => RPIPE_noblock_obuf_3_2_836_inst_req_0); -- 
    outputPort_2_Daemon_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(91) & outputPort_2_Daemon_CP_1176_elements(96);
      gj_outputPort_2_Daemon_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	95 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_3_2_836_update_start_
      -- CP-element group 94: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_3_2_836_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_3_2_836_Update/cr
      -- 
    cr_1379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(94), ack => RPIPE_noblock_obuf_3_2_836_inst_req_1); -- 
    outputPort_2_Daemon_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(92) & outputPort_2_Daemon_CP_1176_elements(95);
      gj_outputPort_2_Daemon_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	94 
    -- CP-element group 95:  members (4) 
      -- CP-element group 95: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_3_2_836_sample_completed__ps
      -- CP-element group 95: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_3_2_836_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_3_2_836_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_3_2_836_Sample/ra
      -- 
    ra_1375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_2_836_inst_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(95)); -- 
    -- CP-element group 96:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	93 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_3_2_836_update_completed__ps
      -- CP-element group 96: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_3_2_836_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_3_2_836_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_3_2_836_Update/ca
      -- 
    ca_1380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_2_836_inst_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(96)); -- 
    -- CP-element group 97:  join  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	9 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	12 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	11 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_837_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	9 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	155 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	13 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_837_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(155);
      gj_outputPort_2_Daemon_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	11 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_837_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(99) <= outputPort_2_Daemon_CP_1176_elements(11);
    -- CP-element group 100:  join  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	12 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_837_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(100) is bound as output of CP function.
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	13 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_837_update_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(101) <= outputPort_2_Daemon_CP_1176_elements(13);
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	154 
    -- CP-element group 102: 	14 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_837_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_837_update_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(102) is bound as output of CP function.
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	7 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_837_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(103) <= outputPort_2_Daemon_CP_1176_elements(7);
    -- CP-element group 104:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_837_loopback_sample_req
      -- CP-element group 104: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_837_loopback_sample_req_ps
      -- 
    phi_stmt_837_loopback_sample_req_1391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_837_loopback_sample_req_1391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(104), ack => phi_stmt_837_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(104) is bound as output of CP function.
    -- CP-element group 105:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	8 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_837_entry_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(105) <= outputPort_2_Daemon_CP_1176_elements(8);
    -- CP-element group 106:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_837_entry_sample_req
      -- CP-element group 106: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_837_entry_sample_req_ps
      -- 
    phi_stmt_837_entry_sample_req_1394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_837_entry_sample_req_1394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(106), ack => phi_stmt_837_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_837_phi_mux_ack
      -- CP-element group 107: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_837_phi_mux_ack_ps
      -- 
    phi_stmt_837_phi_mux_ack_1397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_837_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(107)); -- 
    -- CP-element group 108:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_839_sample_start__ps
      -- CP-element group 108: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_839_sample_completed__ps
      -- CP-element group 108: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_839_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_839_sample_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(108) is bound as output of CP function.
    -- CP-element group 109:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_839_update_start__ps
      -- CP-element group 109: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_839_update_start_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	111 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_839_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(110) <= outputPort_2_Daemon_CP_1176_elements(111);
    -- CP-element group 111:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	110 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_33_839_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(111) is a control-delay.
    cp_element_111_delay: control_delay_element  generic map(name => " 111_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_1176_elements(109), ack => outputPort_2_Daemon_CP_1176_elements(111), clk => clk, reset =>reset);
    -- CP-element group 112:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_4_2_841_sample_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(112) is bound as output of CP function.
    -- CP-element group 113:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_4_2_841_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(113) is bound as output of CP function.
    -- CP-element group 114:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: marked-predecessors 
    -- CP-element group 114: 	117 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_4_2_841_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_4_2_841_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_4_2_841_Sample/rr
      -- 
    rr_1418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(114), ack => RPIPE_noblock_obuf_4_2_841_inst_req_0); -- 
    outputPort_2_Daemon_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(112) & outputPort_2_Daemon_CP_1176_elements(117);
      gj_outputPort_2_Daemon_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	116 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_4_2_841_update_start_
      -- CP-element group 115: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_4_2_841_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_4_2_841_Update/cr
      -- 
    cr_1423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(115), ack => RPIPE_noblock_obuf_4_2_841_inst_req_1); -- 
    outputPort_2_Daemon_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(113) & outputPort_2_Daemon_CP_1176_elements(116);
      gj_outputPort_2_Daemon_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	115 
    -- CP-element group 116:  members (4) 
      -- CP-element group 116: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_4_2_841_sample_completed__ps
      -- CP-element group 116: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_4_2_841_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_4_2_841_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_4_2_841_Sample/ra
      -- 
    ra_1419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_2_841_inst_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(116)); -- 
    -- CP-element group 117:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: marked-successors 
    -- CP-element group 117: 	114 
    -- CP-element group 117:  members (4) 
      -- CP-element group 117: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_4_2_841_update_completed__ps
      -- CP-element group 117: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_4_2_841_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_4_2_841_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/RPIPE_noblock_obuf_4_2_841_Update/ca
      -- 
    ca_1424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_2_841_inst_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(117)); -- 
    -- CP-element group 118:  join  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	9 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	12 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	11 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_842_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  join  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	9 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	155 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	13 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_842_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(155);
      gj_outputPort_2_Daemon_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	11 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_842_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(120) <= outputPort_2_Daemon_CP_1176_elements(11);
    -- CP-element group 121:  join  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	12 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_842_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(121) is bound as output of CP function.
    -- CP-element group 122:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	13 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_842_update_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(122) <= outputPort_2_Daemon_CP_1176_elements(13);
    -- CP-element group 123:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	154 
    -- CP-element group 123: 	14 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_842_update_completed__ps
      -- CP-element group 123: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_842_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(123) is bound as output of CP function.
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	7 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_842_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(124) <= outputPort_2_Daemon_CP_1176_elements(7);
    -- CP-element group 125:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_842_loopback_sample_req_ps
      -- CP-element group 125: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_842_loopback_sample_req
      -- 
    phi_stmt_842_loopback_sample_req_1435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_842_loopback_sample_req_1435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(125), ack => phi_stmt_842_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(125) is bound as output of CP function.
    -- CP-element group 126:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	8 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_842_entry_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(126) <= outputPort_2_Daemon_CP_1176_elements(8);
    -- CP-element group 127:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_842_entry_sample_req_ps
      -- CP-element group 127: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_842_entry_sample_req
      -- 
    phi_stmt_842_entry_sample_req_1438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_842_entry_sample_req_1438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(127), ack => phi_stmt_842_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(127) is bound as output of CP function.
    -- CP-element group 128:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_842_phi_mux_ack
      -- CP-element group 128: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_842_phi_mux_ack_ps
      -- 
    phi_stmt_842_phi_mux_ack_1441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_842_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(128)); -- 
    -- CP-element group 129:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (4) 
      -- CP-element group 129: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_3_844_sample_start_
      -- CP-element group 129: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_3_844_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_3_844_sample_completed__ps
      -- CP-element group 129: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_3_844_sample_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(129) is bound as output of CP function.
    -- CP-element group 130:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (2) 
      -- CP-element group 130: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_3_844_update_start_
      -- CP-element group 130: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_3_844_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(130) is bound as output of CP function.
    -- CP-element group 131:  join  transition  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	132 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_3_844_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(131) <= outputPort_2_Daemon_CP_1176_elements(132);
    -- CP-element group 132:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	131 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ZERO_3_844_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(132) is a control-delay.
    cp_element_132_delay: control_delay_element  generic map(name => " 132_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_1176_elements(130), ack => outputPort_2_Daemon_CP_1176_elements(132), clk => clk, reset =>reset);
    -- CP-element group 133:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	135 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_active_packet_845_Sample/req
      -- CP-element group 133: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_active_packet_845_sample_start__ps
      -- CP-element group 133: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_active_packet_845_Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_active_packet_845_sample_start_
      -- 
    req_1462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(133), ack => next_active_packet_909_845_buf_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(133) is bound as output of CP function.
    -- CP-element group 134:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_active_packet_845_Update/req
      -- CP-element group 134: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_active_packet_845_update_start__ps
      -- CP-element group 134: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_active_packet_845_Update/$entry
      -- CP-element group 134: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_active_packet_845_update_start_
      -- 
    req_1467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(134), ack => next_active_packet_909_845_buf_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(134) is bound as output of CP function.
    -- CP-element group 135:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	133 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (4) 
      -- CP-element group 135: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_active_packet_845_Sample/ack
      -- CP-element group 135: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_active_packet_845_sample_completed__ps
      -- CP-element group 135: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_active_packet_845_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_active_packet_845_sample_completed_
      -- 
    ack_1463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_909_845_buf_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(135)); -- 
    -- CP-element group 136:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (4) 
      -- CP-element group 136: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_active_packet_845_update_completed__ps
      -- CP-element group 136: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_active_packet_845_Update/ack
      -- CP-element group 136: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_active_packet_845_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_active_packet_845_update_completed_
      -- 
    ack_1468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_909_845_buf_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(136)); -- 
    -- CP-element group 137:  join  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	9 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	12 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	11 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_846_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  join  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	9 
    -- CP-element group 138: marked-predecessors 
    -- CP-element group 138: 	155 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	13 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_846_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(155);
      gj_outputPort_2_Daemon_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 139:  join  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	12 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_846_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(139) is bound as output of CP function.
    -- CP-element group 140:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	154 
    -- CP-element group 140: 	14 
    -- CP-element group 140:  members (2) 
      -- CP-element group 140: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_846_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_846_update_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(140) is bound as output of CP function.
    -- CP-element group 141:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	7 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_846_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(141) <= outputPort_2_Daemon_CP_1176_elements(7);
    -- CP-element group 142:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_846_loopback_sample_req
      -- CP-element group 142: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_846_loopback_sample_req_ps
      -- 
    phi_stmt_846_loopback_sample_req_1479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_846_loopback_sample_req_1479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(142), ack => phi_stmt_846_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(142) is bound as output of CP function.
    -- CP-element group 143:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	8 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_846_entry_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(143) <= outputPort_2_Daemon_CP_1176_elements(8);
    -- CP-element group 144:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_846_entry_sample_req
      -- CP-element group 144: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_846_entry_sample_req_ps
      -- 
    phi_stmt_846_entry_sample_req_1482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_846_entry_sample_req_1482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(144), ack => phi_stmt_846_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_846_phi_mux_ack
      -- CP-element group 145: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/phi_stmt_846_phi_mux_ack_ps
      -- 
    phi_stmt_846_phi_mux_ack_1485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_846_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(145)); -- 
    -- CP-element group 146:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (4) 
      -- CP-element group 146: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ONE_3_848_sample_completed_
      -- CP-element group 146: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ONE_3_848_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ONE_3_848_sample_start__ps
      -- CP-element group 146: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ONE_3_848_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(146) is bound as output of CP function.
    -- CP-element group 147:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (2) 
      -- CP-element group 147: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ONE_3_848_update_start_
      -- CP-element group 147: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ONE_3_848_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(147) is bound as output of CP function.
    -- CP-element group 148:  join  transition  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	149 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (1) 
      -- CP-element group 148: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ONE_3_848_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(148) <= outputPort_2_Daemon_CP_1176_elements(149);
    -- CP-element group 149:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	148 
    -- CP-element group 149:  members (1) 
      -- CP-element group 149: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_ONE_3_848_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(149) is a control-delay.
    cp_element_149_delay: control_delay_element  generic map(name => " 149_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_1176_elements(147), ack => outputPort_2_Daemon_CP_1176_elements(149), clk => clk, reset =>reset);
    -- CP-element group 150:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (4) 
      -- CP-element group 150: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_pkt_priority_849_Sample/req
      -- CP-element group 150: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_pkt_priority_849_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_pkt_priority_849_sample_start__ps
      -- CP-element group 150: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_pkt_priority_849_sample_start_
      -- 
    req_1506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(150), ack => next_pkt_priority_909_849_buf_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(150) is bound as output of CP function.
    -- CP-element group 151:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (4) 
      -- CP-element group 151: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_pkt_priority_849_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_pkt_priority_849_Update/req
      -- CP-element group 151: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_pkt_priority_849_update_start_
      -- CP-element group 151: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_pkt_priority_849_update_start__ps
      -- 
    req_1511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(151), ack => next_pkt_priority_909_849_buf_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(151) is bound as output of CP function.
    -- CP-element group 152:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (4) 
      -- CP-element group 152: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_pkt_priority_849_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_pkt_priority_849_Sample/ack
      -- CP-element group 152: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_pkt_priority_849_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_pkt_priority_849_sample_completed__ps
      -- 
    ack_1507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pkt_priority_909_849_buf_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(152)); -- 
    -- CP-element group 153:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (4) 
      -- CP-element group 153: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_pkt_priority_849_Update/ack
      -- CP-element group 153: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_pkt_priority_849_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_pkt_priority_849_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/R_next_pkt_priority_849_update_completed__ps
      -- 
    ack_1512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pkt_priority_909_849_buf_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	140 
    -- CP-element group 154: 	20 
    -- CP-element group 154: 	39 
    -- CP-element group 154: 	60 
    -- CP-element group 154: 	81 
    -- CP-element group 154: 	102 
    -- CP-element group 154: 	123 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/WPIPE_out_data_2_1036_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/WPIPE_out_data_2_1036_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/WPIPE_out_data_2_1036_Sample/req
      -- 
    req_1521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(154), ack => WPIPE_out_data_2_1036_inst_req_0); -- 
    outputPort_2_Daemon_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(140) & outputPort_2_Daemon_CP_1176_elements(20) & outputPort_2_Daemon_CP_1176_elements(39) & outputPort_2_Daemon_CP_1176_elements(60) & outputPort_2_Daemon_CP_1176_elements(81) & outputPort_2_Daemon_CP_1176_elements(102) & outputPort_2_Daemon_CP_1176_elements(123) & outputPort_2_Daemon_CP_1176_elements(156);
      gj_outputPort_2_Daemon_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	138 
    -- CP-element group 155: 	16 
    -- CP-element group 155: 	35 
    -- CP-element group 155: 	56 
    -- CP-element group 155: 	77 
    -- CP-element group 155: 	98 
    -- CP-element group 155: 	119 
    -- CP-element group 155:  members (6) 
      -- CP-element group 155: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/WPIPE_out_data_2_1036_Sample/ack
      -- CP-element group 155: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/WPIPE_out_data_2_1036_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/WPIPE_out_data_2_1036_update_start_
      -- CP-element group 155: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/WPIPE_out_data_2_1036_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/WPIPE_out_data_2_1036_Update/req
      -- CP-element group 155: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/WPIPE_out_data_2_1036_Sample/$exit
      -- 
    ack_1522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_2_1036_inst_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(155)); -- 
    req_1526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(155), ack => WPIPE_out_data_2_1036_inst_req_1); -- 
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	154 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/WPIPE_out_data_2_1036_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/WPIPE_out_data_2_1036_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/WPIPE_out_data_2_1036_Update/ack
      -- 
    ack_1527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_2_1036_inst_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(156)); -- 
    -- CP-element group 157:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	9 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	10 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(157) is a control-delay.
    cp_element_157_delay: control_delay_element  generic map(name => " 157_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_1176_elements(9), ack => outputPort_2_Daemon_CP_1176_elements(157), clk => clk, reset =>reset);
    -- CP-element group 158:  join  transition  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: 	12 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	6 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_815/do_while_stmt_816/do_while_stmt_816_loop_body/$exit
      -- 
    outputPort_2_Daemon_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(156) & outputPort_2_Daemon_CP_1176_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	5 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (2) 
      -- CP-element group 159: 	 branch_block_stmt_815/do_while_stmt_816/loop_exit/$exit
      -- CP-element group 159: 	 branch_block_stmt_815/do_while_stmt_816/loop_exit/ack
      -- 
    ack_1532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_816_branch_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	5 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (2) 
      -- CP-element group 160: 	 branch_block_stmt_815/do_while_stmt_816/loop_taken/ack
      -- CP-element group 160: 	 branch_block_stmt_815/do_while_stmt_816/loop_taken/$exit
      -- 
    ack_1536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_816_branch_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(160)); -- 
    -- CP-element group 161:  transition  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	3 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	1 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_815/do_while_stmt_816/$exit
      -- 
    outputPort_2_Daemon_CP_1176_elements(161) <= outputPort_2_Daemon_CP_1176_elements(3);
    outputPort_2_Daemon_do_while_stmt_816_terminator_1537: loop_terminator -- 
      generic map (name => " outputPort_2_Daemon_do_while_stmt_816_terminator_1537", max_iterations_in_flight =>7) 
      port map(loop_body_exit => outputPort_2_Daemon_CP_1176_elements(6),loop_continue => outputPort_2_Daemon_CP_1176_elements(160),loop_terminate => outputPort_2_Daemon_CP_1176_elements(159),loop_back => outputPort_2_Daemon_CP_1176_elements(4),loop_exit => outputPort_2_Daemon_CP_1176_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_818_phi_seq_1249_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_1176_elements(23);
      outputPort_2_Daemon_CP_1176_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(26);
      outputPort_2_Daemon_CP_1176_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(28);
      outputPort_2_Daemon_CP_1176_elements(24) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_1176_elements(21);
      outputPort_2_Daemon_CP_1176_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(32);
      outputPort_2_Daemon_CP_1176_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(33);
      outputPort_2_Daemon_CP_1176_elements(22) <= phi_mux_reqs(1);
      phi_stmt_818_phi_seq_1249 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_818_phi_seq_1249") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_1176_elements(17), 
          phi_sample_ack => outputPort_2_Daemon_CP_1176_elements(18), 
          phi_update_req => outputPort_2_Daemon_CP_1176_elements(19), 
          phi_update_ack => outputPort_2_Daemon_CP_1176_elements(20), 
          phi_mux_ack => outputPort_2_Daemon_CP_1176_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_822_phi_seq_1293_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_1176_elements(42);
      outputPort_2_Daemon_CP_1176_elements(45)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(45);
      outputPort_2_Daemon_CP_1176_elements(46)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(47);
      outputPort_2_Daemon_CP_1176_elements(43) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_1176_elements(40);
      outputPort_2_Daemon_CP_1176_elements(49)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(53);
      outputPort_2_Daemon_CP_1176_elements(50)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(54);
      outputPort_2_Daemon_CP_1176_elements(41) <= phi_mux_reqs(1);
      phi_stmt_822_phi_seq_1293 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_822_phi_seq_1293") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_1176_elements(36), 
          phi_sample_ack => outputPort_2_Daemon_CP_1176_elements(37), 
          phi_update_req => outputPort_2_Daemon_CP_1176_elements(38), 
          phi_update_ack => outputPort_2_Daemon_CP_1176_elements(39), 
          phi_mux_ack => outputPort_2_Daemon_CP_1176_elements(44), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_827_phi_seq_1337_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_1176_elements(63);
      outputPort_2_Daemon_CP_1176_elements(66)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(66);
      outputPort_2_Daemon_CP_1176_elements(67)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(68);
      outputPort_2_Daemon_CP_1176_elements(64) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_1176_elements(61);
      outputPort_2_Daemon_CP_1176_elements(70)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(74);
      outputPort_2_Daemon_CP_1176_elements(71)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(75);
      outputPort_2_Daemon_CP_1176_elements(62) <= phi_mux_reqs(1);
      phi_stmt_827_phi_seq_1337 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_827_phi_seq_1337") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_1176_elements(57), 
          phi_sample_ack => outputPort_2_Daemon_CP_1176_elements(58), 
          phi_update_req => outputPort_2_Daemon_CP_1176_elements(59), 
          phi_update_ack => outputPort_2_Daemon_CP_1176_elements(60), 
          phi_mux_ack => outputPort_2_Daemon_CP_1176_elements(65), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_832_phi_seq_1381_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_1176_elements(84);
      outputPort_2_Daemon_CP_1176_elements(87)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(87);
      outputPort_2_Daemon_CP_1176_elements(88)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(89);
      outputPort_2_Daemon_CP_1176_elements(85) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_1176_elements(82);
      outputPort_2_Daemon_CP_1176_elements(91)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(95);
      outputPort_2_Daemon_CP_1176_elements(92)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(96);
      outputPort_2_Daemon_CP_1176_elements(83) <= phi_mux_reqs(1);
      phi_stmt_832_phi_seq_1381 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_832_phi_seq_1381") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_1176_elements(78), 
          phi_sample_ack => outputPort_2_Daemon_CP_1176_elements(79), 
          phi_update_req => outputPort_2_Daemon_CP_1176_elements(80), 
          phi_update_ack => outputPort_2_Daemon_CP_1176_elements(81), 
          phi_mux_ack => outputPort_2_Daemon_CP_1176_elements(86), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_837_phi_seq_1425_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_1176_elements(105);
      outputPort_2_Daemon_CP_1176_elements(108)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(108);
      outputPort_2_Daemon_CP_1176_elements(109)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(110);
      outputPort_2_Daemon_CP_1176_elements(106) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_1176_elements(103);
      outputPort_2_Daemon_CP_1176_elements(112)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(116);
      outputPort_2_Daemon_CP_1176_elements(113)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(117);
      outputPort_2_Daemon_CP_1176_elements(104) <= phi_mux_reqs(1);
      phi_stmt_837_phi_seq_1425 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_837_phi_seq_1425") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_1176_elements(99), 
          phi_sample_ack => outputPort_2_Daemon_CP_1176_elements(100), 
          phi_update_req => outputPort_2_Daemon_CP_1176_elements(101), 
          phi_update_ack => outputPort_2_Daemon_CP_1176_elements(102), 
          phi_mux_ack => outputPort_2_Daemon_CP_1176_elements(107), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_842_phi_seq_1469_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_1176_elements(126);
      outputPort_2_Daemon_CP_1176_elements(129)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(129);
      outputPort_2_Daemon_CP_1176_elements(130)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(131);
      outputPort_2_Daemon_CP_1176_elements(127) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_1176_elements(124);
      outputPort_2_Daemon_CP_1176_elements(133)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(135);
      outputPort_2_Daemon_CP_1176_elements(134)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(136);
      outputPort_2_Daemon_CP_1176_elements(125) <= phi_mux_reqs(1);
      phi_stmt_842_phi_seq_1469 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_842_phi_seq_1469") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_1176_elements(120), 
          phi_sample_ack => outputPort_2_Daemon_CP_1176_elements(121), 
          phi_update_req => outputPort_2_Daemon_CP_1176_elements(122), 
          phi_update_ack => outputPort_2_Daemon_CP_1176_elements(123), 
          phi_mux_ack => outputPort_2_Daemon_CP_1176_elements(128), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_846_phi_seq_1513_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_1176_elements(143);
      outputPort_2_Daemon_CP_1176_elements(146)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(146);
      outputPort_2_Daemon_CP_1176_elements(147)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(148);
      outputPort_2_Daemon_CP_1176_elements(144) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_1176_elements(141);
      outputPort_2_Daemon_CP_1176_elements(150)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(152);
      outputPort_2_Daemon_CP_1176_elements(151)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(153);
      outputPort_2_Daemon_CP_1176_elements(142) <= phi_mux_reqs(1);
      phi_stmt_846_phi_seq_1513 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_846_phi_seq_1513") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_1176_elements(11), 
          phi_sample_ack => outputPort_2_Daemon_CP_1176_elements(139), 
          phi_update_req => outputPort_2_Daemon_CP_1176_elements(13), 
          phi_update_ack => outputPort_2_Daemon_CP_1176_elements(140), 
          phi_mux_ack => outputPort_2_Daemon_CP_1176_elements(145), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1201_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= outputPort_2_Daemon_CP_1176_elements(7);
        preds(1)  <= outputPort_2_Daemon_CP_1176_elements(8);
        entry_tmerge_1201 : transition_merge -- 
          generic map(name => " entry_tmerge_1201")
          port map (preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u3_u1_1009_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1015_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1022_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1028_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_874_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_880_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_887_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_893_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_935_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_943_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_951_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_959_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_976_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_983_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_991_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_998_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_916_wire : std_logic_vector(0 downto 0);
    signal MUX_1002_wire : std_logic_vector(31 downto 0);
    signal MUX_1012_wire : std_logic_vector(0 downto 0);
    signal MUX_1018_wire : std_logic_vector(0 downto 0);
    signal MUX_1025_wire : std_logic_vector(0 downto 0);
    signal MUX_1031_wire : std_logic_vector(0 downto 0);
    signal MUX_877_wire : std_logic_vector(0 downto 0);
    signal MUX_883_wire : std_logic_vector(0 downto 0);
    signal MUX_890_wire : std_logic_vector(0 downto 0);
    signal MUX_896_wire : std_logic_vector(0 downto 0);
    signal MUX_927_wire : std_logic_vector(7 downto 0);
    signal MUX_980_wire : std_logic_vector(31 downto 0);
    signal MUX_987_wire : std_logic_vector(31 downto 0);
    signal MUX_995_wire : std_logic_vector(31 downto 0);
    signal NEQ_u3_u1_913_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_932_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_940_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_948_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_956_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1019_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1032_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_884_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_897_wire : std_logic_vector(0 downto 0);
    signal OR_u32_u32_1003_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_988_wire : std_logic_vector(31 downto 0);
    signal RPIPE_noblock_obuf_1_2_826_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_2_2_831_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_3_2_836_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_4_2_841_wire : std_logic_vector(32 downto 0);
    signal R_ONE_3_848_wire_constant : std_logic_vector(2 downto 0);
    signal R_ZERO_33_824_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_829_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_834_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_839_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_3_844_wire_constant : std_logic_vector(2 downto 0);
    signal R_ZERO_8_820_wire_constant : std_logic_vector(7 downto 0);
    signal SUB_u8_u8_925_wire : std_logic_vector(7 downto 0);
    signal active_packet_842 : std_logic_vector(2 downto 0);
    signal data_to_out_1005 : std_logic_vector(31 downto 0);
    signal down_counter_818 : std_logic_vector(7 downto 0);
    signal konst_1001_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1008_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1011_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1014_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1017_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1021_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1024_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1027_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1030_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1040_wire_constant : std_logic_vector(0 downto 0);
    signal konst_853_wire_constant : std_logic_vector(32 downto 0);
    signal konst_858_wire_constant : std_logic_vector(32 downto 0);
    signal konst_863_wire_constant : std_logic_vector(32 downto 0);
    signal konst_868_wire_constant : std_logic_vector(32 downto 0);
    signal konst_873_wire_constant : std_logic_vector(2 downto 0);
    signal konst_876_wire_constant : std_logic_vector(0 downto 0);
    signal konst_879_wire_constant : std_logic_vector(2 downto 0);
    signal konst_882_wire_constant : std_logic_vector(0 downto 0);
    signal konst_886_wire_constant : std_logic_vector(2 downto 0);
    signal konst_889_wire_constant : std_logic_vector(0 downto 0);
    signal konst_892_wire_constant : std_logic_vector(2 downto 0);
    signal konst_895_wire_constant : std_logic_vector(0 downto 0);
    signal konst_912_wire_constant : std_logic_vector(2 downto 0);
    signal konst_915_wire_constant : std_logic_vector(7 downto 0);
    signal konst_921_wire_constant : std_logic_vector(7 downto 0);
    signal konst_924_wire_constant : std_logic_vector(7 downto 0);
    signal konst_934_wire_constant : std_logic_vector(2 downto 0);
    signal konst_942_wire_constant : std_logic_vector(2 downto 0);
    signal konst_950_wire_constant : std_logic_vector(2 downto 0);
    signal konst_958_wire_constant : std_logic_vector(2 downto 0);
    signal konst_975_wire_constant : std_logic_vector(2 downto 0);
    signal konst_979_wire_constant : std_logic_vector(31 downto 0);
    signal konst_982_wire_constant : std_logic_vector(2 downto 0);
    signal konst_986_wire_constant : std_logic_vector(31 downto 0);
    signal konst_990_wire_constant : std_logic_vector(2 downto 0);
    signal konst_994_wire_constant : std_logic_vector(31 downto 0);
    signal konst_997_wire_constant : std_logic_vector(2 downto 0);
    signal next_active_packet_909 : std_logic_vector(2 downto 0);
    signal next_active_packet_909_845_buffered : std_logic_vector(2 downto 0);
    signal next_down_counter_929 : std_logic_vector(7 downto 0);
    signal next_down_counter_929_821_buffered : std_logic_vector(7 downto 0);
    signal next_pkt_priority_909 : std_logic_vector(2 downto 0);
    signal next_pkt_priority_909_849_buffered : std_logic_vector(2 downto 0);
    signal p1_valid_855 : std_logic_vector(0 downto 0);
    signal p2_valid_860 : std_logic_vector(0 downto 0);
    signal p3_valid_865 : std_logic_vector(0 downto 0);
    signal p4_valid_870 : std_logic_vector(0 downto 0);
    signal pkt_1_e_word_822 : std_logic_vector(32 downto 0);
    signal pkt_2_e_word_827 : std_logic_vector(32 downto 0);
    signal pkt_3_e_word_832 : std_logic_vector(32 downto 0);
    signal pkt_4_e_word_837 : std_logic_vector(32 downto 0);
    signal pkt_priority_846 : std_logic_vector(2 downto 0);
    signal read_from_1_937 : std_logic_vector(0 downto 0);
    signal read_from_2_945 : std_logic_vector(0 downto 0);
    signal read_from_3_953 : std_logic_vector(0 downto 0);
    signal read_from_4_961 : std_logic_vector(0 downto 0);
    signal send_flag_1034 : std_logic_vector(0 downto 0);
    signal slice_1000_wire : std_logic_vector(31 downto 0);
    signal slice_978_wire : std_logic_vector(31 downto 0);
    signal slice_985_wire : std_logic_vector(31 downto 0);
    signal slice_993_wire : std_logic_vector(31 downto 0);
    signal started_new_packet_918 : std_logic_vector(0 downto 0);
    signal valid_active_pkt_word_read_899 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_ONE_3_848_wire_constant <= "001";
    R_ZERO_33_824_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_829_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_834_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_839_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_3_844_wire_constant <= "000";
    R_ZERO_8_820_wire_constant <= "00000000";
    konst_1001_wire_constant <= "00000000000000000000000000000000";
    konst_1008_wire_constant <= "001";
    konst_1011_wire_constant <= "0";
    konst_1014_wire_constant <= "010";
    konst_1017_wire_constant <= "0";
    konst_1021_wire_constant <= "011";
    konst_1024_wire_constant <= "0";
    konst_1027_wire_constant <= "100";
    konst_1030_wire_constant <= "0";
    konst_1040_wire_constant <= "1";
    konst_853_wire_constant <= "000000000000000000000000000100000";
    konst_858_wire_constant <= "000000000000000000000000000100000";
    konst_863_wire_constant <= "000000000000000000000000000100000";
    konst_868_wire_constant <= "000000000000000000000000000100000";
    konst_873_wire_constant <= "001";
    konst_876_wire_constant <= "0";
    konst_879_wire_constant <= "010";
    konst_882_wire_constant <= "0";
    konst_886_wire_constant <= "011";
    konst_889_wire_constant <= "0";
    konst_892_wire_constant <= "100";
    konst_895_wire_constant <= "0";
    konst_912_wire_constant <= "000";
    konst_915_wire_constant <= "00000000";
    konst_921_wire_constant <= "00111111";
    konst_924_wire_constant <= "00000001";
    konst_934_wire_constant <= "001";
    konst_942_wire_constant <= "010";
    konst_950_wire_constant <= "011";
    konst_958_wire_constant <= "100";
    konst_975_wire_constant <= "001";
    konst_979_wire_constant <= "00000000000000000000000000000000";
    konst_982_wire_constant <= "010";
    konst_986_wire_constant <= "00000000000000000000000000000000";
    konst_990_wire_constant <= "011";
    konst_994_wire_constant <= "00000000000000000000000000000000";
    konst_997_wire_constant <= "100";
    phi_stmt_818: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_8_820_wire_constant & next_down_counter_929_821_buffered;
      req <= phi_stmt_818_req_0 & phi_stmt_818_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_818",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_818_ack_0,
          idata => idata,
          odata => down_counter_818,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_818
    phi_stmt_822: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_824_wire_constant & RPIPE_noblock_obuf_1_2_826_wire;
      req <= phi_stmt_822_req_0 & phi_stmt_822_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_822",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_822_ack_0,
          idata => idata,
          odata => pkt_1_e_word_822,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_822
    phi_stmt_827: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_829_wire_constant & RPIPE_noblock_obuf_2_2_831_wire;
      req <= phi_stmt_827_req_0 & phi_stmt_827_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_827",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_827_ack_0,
          idata => idata,
          odata => pkt_2_e_word_827,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_827
    phi_stmt_832: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_834_wire_constant & RPIPE_noblock_obuf_3_2_836_wire;
      req <= phi_stmt_832_req_0 & phi_stmt_832_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_832",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_832_ack_0,
          idata => idata,
          odata => pkt_3_e_word_832,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_832
    phi_stmt_837: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_839_wire_constant & RPIPE_noblock_obuf_4_2_841_wire;
      req <= phi_stmt_837_req_0 & phi_stmt_837_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_837",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_837_ack_0,
          idata => idata,
          odata => pkt_4_e_word_837,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_837
    phi_stmt_842: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_3_844_wire_constant & next_active_packet_909_845_buffered;
      req <= phi_stmt_842_req_0 & phi_stmt_842_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_842",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_842_ack_0,
          idata => idata,
          odata => active_packet_842,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_842
    phi_stmt_846: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ONE_3_848_wire_constant & next_pkt_priority_909_849_buffered;
      req <= phi_stmt_846_req_0 & phi_stmt_846_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_846",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_846_ack_0,
          idata => idata,
          odata => pkt_priority_846,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_846
    -- flow-through select operator MUX_1002_inst
    MUX_1002_wire <= slice_1000_wire when (EQ_u3_u1_998_wire(0) /=  '0') else konst_1001_wire_constant;
    -- flow-through select operator MUX_1012_inst
    MUX_1012_wire <= p1_valid_855 when (EQ_u3_u1_1009_wire(0) /=  '0') else konst_1011_wire_constant;
    -- flow-through select operator MUX_1018_inst
    MUX_1018_wire <= p2_valid_860 when (EQ_u3_u1_1015_wire(0) /=  '0') else konst_1017_wire_constant;
    -- flow-through select operator MUX_1025_inst
    MUX_1025_wire <= p3_valid_865 when (EQ_u3_u1_1022_wire(0) /=  '0') else konst_1024_wire_constant;
    -- flow-through select operator MUX_1031_inst
    MUX_1031_wire <= p4_valid_870 when (EQ_u3_u1_1028_wire(0) /=  '0') else konst_1030_wire_constant;
    -- flow-through select operator MUX_877_inst
    MUX_877_wire <= p1_valid_855 when (EQ_u3_u1_874_wire(0) /=  '0') else konst_876_wire_constant;
    -- flow-through select operator MUX_883_inst
    MUX_883_wire <= p2_valid_860 when (EQ_u3_u1_880_wire(0) /=  '0') else konst_882_wire_constant;
    -- flow-through select operator MUX_890_inst
    MUX_890_wire <= p3_valid_865 when (EQ_u3_u1_887_wire(0) /=  '0') else konst_889_wire_constant;
    -- flow-through select operator MUX_896_inst
    MUX_896_wire <= p4_valid_870 when (EQ_u3_u1_893_wire(0) /=  '0') else konst_895_wire_constant;
    -- flow-through select operator MUX_927_inst
    MUX_927_wire <= SUB_u8_u8_925_wire when (valid_active_pkt_word_read_899(0) /=  '0') else down_counter_818;
    -- flow-through select operator MUX_928_inst
    next_down_counter_929 <= konst_921_wire_constant when (started_new_packet_918(0) /=  '0') else MUX_927_wire;
    -- flow-through select operator MUX_980_inst
    MUX_980_wire <= slice_978_wire when (EQ_u3_u1_976_wire(0) /=  '0') else konst_979_wire_constant;
    -- flow-through select operator MUX_987_inst
    MUX_987_wire <= slice_985_wire when (EQ_u3_u1_983_wire(0) /=  '0') else konst_986_wire_constant;
    -- flow-through select operator MUX_995_inst
    MUX_995_wire <= slice_993_wire when (EQ_u3_u1_991_wire(0) /=  '0') else konst_994_wire_constant;
    -- flow-through slice operator slice_1000_inst
    slice_1000_wire <= pkt_4_e_word_837(31 downto 0);
    -- flow-through slice operator slice_978_inst
    slice_978_wire <= pkt_1_e_word_822(31 downto 0);
    -- flow-through slice operator slice_985_inst
    slice_985_wire <= pkt_2_e_word_827(31 downto 0);
    -- flow-through slice operator slice_993_inst
    slice_993_wire <= pkt_3_e_word_832(31 downto 0);
    next_active_packet_909_845_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_active_packet_909_845_buf_req_0;
      next_active_packet_909_845_buf_ack_0<= wack(0);
      rreq(0) <= next_active_packet_909_845_buf_req_1;
      next_active_packet_909_845_buf_ack_1<= rack(0);
      next_active_packet_909_845_buf : InterlockBuffer generic map ( -- 
        name => "next_active_packet_909_845_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_active_packet_909,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_active_packet_909_845_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_down_counter_929_821_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_down_counter_929_821_buf_req_0;
      next_down_counter_929_821_buf_ack_0<= wack(0);
      rreq(0) <= next_down_counter_929_821_buf_req_1;
      next_down_counter_929_821_buf_ack_1<= rack(0);
      next_down_counter_929_821_buf : InterlockBuffer generic map ( -- 
        name => "next_down_counter_929_821_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_down_counter_929,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_down_counter_929_821_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_pkt_priority_909_849_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_pkt_priority_909_849_buf_req_0;
      next_pkt_priority_909_849_buf_ack_0<= wack(0);
      rreq(0) <= next_pkt_priority_909_849_buf_req_1;
      next_pkt_priority_909_849_buf_ack_1<= rack(0);
      next_pkt_priority_909_849_buf : InterlockBuffer generic map ( -- 
        name => "next_pkt_priority_909_849_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_pkt_priority_909,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_pkt_priority_909_849_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_816_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1040_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_816_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_816_branch_req_0,
          ack0 => do_while_stmt_816_branch_ack_0,
          ack1 => do_while_stmt_816_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator AND_u1_u1_917_inst
    process(NEQ_u3_u1_913_wire, EQ_u8_u1_916_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NEQ_u3_u1_913_wire, EQ_u8_u1_916_wire, tmp_var);
      started_new_packet_918 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_854_inst
    process(pkt_1_e_word_822) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_1_e_word_822, konst_853_wire_constant, tmp_var);
      p1_valid_855 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_859_inst
    process(pkt_2_e_word_827) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_2_e_word_827, konst_858_wire_constant, tmp_var);
      p2_valid_860 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_864_inst
    process(pkt_3_e_word_832) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_3_e_word_832, konst_863_wire_constant, tmp_var);
      p3_valid_865 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_869_inst
    process(pkt_4_e_word_837) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_4_e_word_837, konst_868_wire_constant, tmp_var);
      p4_valid_870 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1009_inst
    process(next_active_packet_909) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_909, konst_1008_wire_constant, tmp_var);
      EQ_u3_u1_1009_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1015_inst
    process(next_active_packet_909) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_909, konst_1014_wire_constant, tmp_var);
      EQ_u3_u1_1015_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1022_inst
    process(next_active_packet_909) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_909, konst_1021_wire_constant, tmp_var);
      EQ_u3_u1_1022_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1028_inst
    process(next_active_packet_909) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_909, konst_1027_wire_constant, tmp_var);
      EQ_u3_u1_1028_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_874_inst
    process(active_packet_842) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_842, konst_873_wire_constant, tmp_var);
      EQ_u3_u1_874_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_880_inst
    process(active_packet_842) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_842, konst_879_wire_constant, tmp_var);
      EQ_u3_u1_880_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_887_inst
    process(active_packet_842) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_842, konst_886_wire_constant, tmp_var);
      EQ_u3_u1_887_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_893_inst
    process(active_packet_842) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_842, konst_892_wire_constant, tmp_var);
      EQ_u3_u1_893_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_935_inst
    process(next_active_packet_909) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_909, konst_934_wire_constant, tmp_var);
      EQ_u3_u1_935_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_943_inst
    process(next_active_packet_909) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_909, konst_942_wire_constant, tmp_var);
      EQ_u3_u1_943_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_951_inst
    process(next_active_packet_909) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_909, konst_950_wire_constant, tmp_var);
      EQ_u3_u1_951_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_959_inst
    process(next_active_packet_909) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_909, konst_958_wire_constant, tmp_var);
      EQ_u3_u1_959_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_976_inst
    process(next_active_packet_909) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_909, konst_975_wire_constant, tmp_var);
      EQ_u3_u1_976_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_983_inst
    process(next_active_packet_909) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_909, konst_982_wire_constant, tmp_var);
      EQ_u3_u1_983_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_991_inst
    process(next_active_packet_909) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_909, konst_990_wire_constant, tmp_var);
      EQ_u3_u1_991_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_998_inst
    process(next_active_packet_909) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_909, konst_997_wire_constant, tmp_var);
      EQ_u3_u1_998_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_916_inst
    process(down_counter_818) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(down_counter_818, konst_915_wire_constant, tmp_var);
      EQ_u8_u1_916_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u3_u1_913_inst
    process(next_active_packet_909) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(next_active_packet_909, konst_912_wire_constant, tmp_var);
      NEQ_u3_u1_913_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_932_inst
    process(p1_valid_855) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_855, tmp_var);
      NOT_u1_u1_932_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_940_inst
    process(p2_valid_860) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_860, tmp_var);
      NOT_u1_u1_940_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_948_inst
    process(p3_valid_865) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_865, tmp_var);
      NOT_u1_u1_948_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_956_inst
    process(p4_valid_870) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_870, tmp_var);
      NOT_u1_u1_956_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1019_inst
    process(MUX_1012_wire, MUX_1018_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1012_wire, MUX_1018_wire, tmp_var);
      OR_u1_u1_1019_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1032_inst
    process(MUX_1025_wire, MUX_1031_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1025_wire, MUX_1031_wire, tmp_var);
      OR_u1_u1_1032_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1033_inst
    process(OR_u1_u1_1019_wire, OR_u1_u1_1032_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1019_wire, OR_u1_u1_1032_wire, tmp_var);
      send_flag_1034 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_884_inst
    process(MUX_877_wire, MUX_883_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_877_wire, MUX_883_wire, tmp_var);
      OR_u1_u1_884_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_897_inst
    process(MUX_890_wire, MUX_896_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_890_wire, MUX_896_wire, tmp_var);
      OR_u1_u1_897_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_898_inst
    process(OR_u1_u1_884_wire, OR_u1_u1_897_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_884_wire, OR_u1_u1_897_wire, tmp_var);
      valid_active_pkt_word_read_899 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_936_inst
    process(NOT_u1_u1_932_wire, EQ_u3_u1_935_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_932_wire, EQ_u3_u1_935_wire, tmp_var);
      read_from_1_937 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_944_inst
    process(NOT_u1_u1_940_wire, EQ_u3_u1_943_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_940_wire, EQ_u3_u1_943_wire, tmp_var);
      read_from_2_945 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_952_inst
    process(NOT_u1_u1_948_wire, EQ_u3_u1_951_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_948_wire, EQ_u3_u1_951_wire, tmp_var);
      read_from_3_953 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_960_inst
    process(NOT_u1_u1_956_wire, EQ_u3_u1_959_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_956_wire, EQ_u3_u1_959_wire, tmp_var);
      read_from_4_961 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1003_inst
    process(MUX_995_wire, MUX_1002_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_995_wire, MUX_1002_wire, tmp_var);
      OR_u32_u32_1003_wire <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1004_inst
    process(OR_u32_u32_988_wire, OR_u32_u32_1003_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u32_u32_988_wire, OR_u32_u32_1003_wire, tmp_var);
      data_to_out_1005 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_988_inst
    process(MUX_980_wire, MUX_987_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_980_wire, MUX_987_wire, tmp_var);
      OR_u32_u32_988_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u8_u8_925_inst
    process(down_counter_818) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSub_proc(down_counter_818, konst_924_wire_constant, tmp_var);
      SUB_u8_u8_925_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_noblock_obuf_1_2_826_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_1_2_826_inst_req_0;
      RPIPE_noblock_obuf_1_2_826_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_1_2_826_inst_req_1;
      RPIPE_noblock_obuf_1_2_826_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_1_937(0);
      RPIPE_noblock_obuf_1_2_826_wire <= data_out(32 downto 0);
      noblock_obuf_1_2_read_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_2_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_2_read_0: InputPortRevised -- 
        generic map ( name => "noblock_obuf_1_2_read_0", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_1_2_pipe_read_req(0),
          oack => noblock_obuf_1_2_pipe_read_ack(0),
          odata => noblock_obuf_1_2_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_noblock_obuf_2_2_831_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_2_2_831_inst_req_0;
      RPIPE_noblock_obuf_2_2_831_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_2_2_831_inst_req_1;
      RPIPE_noblock_obuf_2_2_831_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_2_945(0);
      RPIPE_noblock_obuf_2_2_831_wire <= data_out(32 downto 0);
      noblock_obuf_2_2_read_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_2_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_2_read_1: InputPortRevised -- 
        generic map ( name => "noblock_obuf_2_2_read_1", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_2_2_pipe_read_req(0),
          oack => noblock_obuf_2_2_pipe_read_ack(0),
          odata => noblock_obuf_2_2_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_noblock_obuf_3_2_836_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_3_2_836_inst_req_0;
      RPIPE_noblock_obuf_3_2_836_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_3_2_836_inst_req_1;
      RPIPE_noblock_obuf_3_2_836_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_3_953(0);
      RPIPE_noblock_obuf_3_2_836_wire <= data_out(32 downto 0);
      noblock_obuf_3_2_read_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_2_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_2_read_2: InputPortRevised -- 
        generic map ( name => "noblock_obuf_3_2_read_2", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_3_2_pipe_read_req(0),
          oack => noblock_obuf_3_2_pipe_read_ack(0),
          odata => noblock_obuf_3_2_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_noblock_obuf_4_2_841_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_4_2_841_inst_req_0;
      RPIPE_noblock_obuf_4_2_841_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_4_2_841_inst_req_1;
      RPIPE_noblock_obuf_4_2_841_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_4_961(0);
      RPIPE_noblock_obuf_4_2_841_wire <= data_out(32 downto 0);
      noblock_obuf_4_2_read_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_2_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_2_read_3: InputPortRevised -- 
        generic map ( name => "noblock_obuf_4_2_read_3", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_4_2_pipe_read_req(0),
          oack => noblock_obuf_4_2_pipe_read_ack(0),
          odata => noblock_obuf_4_2_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_out_data_2_1036_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_out_data_2_1036_inst_req_0;
      WPIPE_out_data_2_1036_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_out_data_2_1036_inst_req_1;
      WPIPE_out_data_2_1036_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_flag_1034(0);
      data_in <= data_to_out_1005;
      out_data_2_write_0_gI: SplitGuardInterface generic map(name => "out_data_2_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      out_data_2_write_0: OutputPortRevised -- 
        generic map ( name => "out_data_2", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => out_data_2_pipe_write_req(0),
          oack => out_data_2_pipe_write_ack(0),
          odata => out_data_2_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    volatile_operator_prioritySelect_2477: prioritySelect_Volatile port map(down_counter => down_counter_818, active_packet => active_packet_842, pkt_priority => pkt_priority_846, p1_valid => p1_valid_855, p2_valid => p2_valid_860, p3_valid => p3_valid_865, p4_valid => p4_valid_870, next_active_packet => next_active_packet_909, next_pkt_priority => next_pkt_priority_909); 
    -- 
  end Block; -- data_path
  -- 
end outputPort_2_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity outputPort_3_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    noblock_obuf_1_3_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_3_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_3_3_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_3_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_4_3_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_3_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_2_3_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_3_pipe_read_data : in   std_logic_vector(32 downto 0);
    out_data_3_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_3_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity outputPort_3_Daemon;
architecture outputPort_3_Daemon_arch of outputPort_3_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal outputPort_3_Daemon_CP_1538_start: Boolean;
  signal outputPort_3_Daemon_CP_1538_symbol: Boolean;
  -- volatile/operator module components. 
  component prioritySelect_Volatile is -- 
    port ( -- 
      down_counter : in  std_logic_vector(7 downto 0);
      active_packet : in  std_logic_vector(2 downto 0);
      pkt_priority : in  std_logic_vector(2 downto 0);
      p1_valid : in  std_logic_vector(0 downto 0);
      p2_valid : in  std_logic_vector(0 downto 0);
      p3_valid : in  std_logic_vector(0 downto 0);
      p4_valid : in  std_logic_vector(0 downto 0);
      next_active_packet : out  std_logic_vector(2 downto 0);
      next_pkt_priority : out  std_logic_vector(2 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal RPIPE_noblock_obuf_3_3_1065_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_3_3_1065_inst_req_0 : boolean;
  signal do_while_stmt_1045_branch_ack_0 : boolean;
  signal next_active_packet_1138_1074_buf_req_0 : boolean;
  signal next_pkt_priority_1138_1078_buf_req_0 : boolean;
  signal next_pkt_priority_1138_1078_buf_req_1 : boolean;
  signal phi_stmt_1071_req_1 : boolean;
  signal next_pkt_priority_1138_1078_buf_ack_0 : boolean;
  signal next_pkt_priority_1138_1078_buf_ack_1 : boolean;
  signal WPIPE_out_data_3_1265_inst_ack_1 : boolean;
  signal RPIPE_noblock_obuf_4_3_1070_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_4_3_1070_inst_ack_0 : boolean;
  signal next_active_packet_1138_1074_buf_ack_1 : boolean;
  signal WPIPE_out_data_3_1265_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_4_3_1070_inst_ack_1 : boolean;
  signal phi_stmt_1066_req_1 : boolean;
  signal next_active_packet_1138_1074_buf_req_1 : boolean;
  signal next_active_packet_1138_1074_buf_ack_0 : boolean;
  signal phi_stmt_1066_req_0 : boolean;
  signal do_while_stmt_1045_branch_ack_1 : boolean;
  signal phi_stmt_1075_req_1 : boolean;
  signal phi_stmt_1075_req_0 : boolean;
  signal RPIPE_noblock_obuf_3_3_1065_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_3_3_1065_inst_ack_1 : boolean;
  signal phi_stmt_1075_ack_0 : boolean;
  signal phi_stmt_1066_ack_0 : boolean;
  signal WPIPE_out_data_3_1265_inst_req_0 : boolean;
  signal WPIPE_out_data_3_1265_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_4_3_1070_inst_req_0 : boolean;
  signal phi_stmt_1071_ack_0 : boolean;
  signal phi_stmt_1071_req_0 : boolean;
  signal do_while_stmt_1045_branch_req_0 : boolean;
  signal phi_stmt_1047_req_1 : boolean;
  signal phi_stmt_1047_req_0 : boolean;
  signal phi_stmt_1047_ack_0 : boolean;
  signal next_down_counter_1158_1050_buf_req_0 : boolean;
  signal next_down_counter_1158_1050_buf_ack_0 : boolean;
  signal next_down_counter_1158_1050_buf_req_1 : boolean;
  signal next_down_counter_1158_1050_buf_ack_1 : boolean;
  signal phi_stmt_1051_req_1 : boolean;
  signal phi_stmt_1051_req_0 : boolean;
  signal phi_stmt_1051_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_3_1055_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_1_3_1055_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_3_1055_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_1_3_1055_inst_ack_1 : boolean;
  signal phi_stmt_1056_req_1 : boolean;
  signal phi_stmt_1056_req_0 : boolean;
  signal phi_stmt_1056_ack_0 : boolean;
  signal RPIPE_noblock_obuf_2_3_1060_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_2_3_1060_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_2_3_1060_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_2_3_1060_inst_ack_1 : boolean;
  signal phi_stmt_1061_req_1 : boolean;
  signal phi_stmt_1061_req_0 : boolean;
  signal phi_stmt_1061_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "outputPort_3_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  outputPort_3_Daemon_CP_1538_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "outputPort_3_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_3_Daemon_CP_1538_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= outputPort_3_Daemon_CP_1538_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_3_Daemon_CP_1538_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  outputPort_3_Daemon_CP_1538: Block -- control-path 
    signal outputPort_3_Daemon_CP_1538_elements: BooleanArray(161 downto 0);
    -- 
  begin -- 
    outputPort_3_Daemon_CP_1538_elements(0) <= outputPort_3_Daemon_CP_1538_start;
    outputPort_3_Daemon_CP_1538_symbol <= outputPort_3_Daemon_CP_1538_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1044/$entry
      -- CP-element group 0: 	 branch_block_stmt_1044/branch_block_stmt_1044__entry__
      -- CP-element group 0: 	 branch_block_stmt_1044/do_while_stmt_1045__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	161 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1044/$exit
      -- CP-element group 1: 	 branch_block_stmt_1044/branch_block_stmt_1044__exit__
      -- CP-element group 1: 	 branch_block_stmt_1044/do_while_stmt_1045__exit__
      -- 
    outputPort_3_Daemon_CP_1538_elements(1) <= outputPort_3_Daemon_CP_1538_elements(161);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1044/do_while_stmt_1045/$entry
      -- CP-element group 2: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045__entry__
      -- 
    outputPort_3_Daemon_CP_1538_elements(2) <= outputPort_3_Daemon_CP_1538_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	161 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045__exit__
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1044/do_while_stmt_1045/loop_back
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	160 
    -- CP-element group 5: 	159 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1044/do_while_stmt_1045/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1044/do_while_stmt_1045/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_1044/do_while_stmt_1045/condition_done
      -- 
    outputPort_3_Daemon_CP_1538_elements(5) <= outputPort_3_Daemon_CP_1538_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	158 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1044/do_while_stmt_1045/loop_body_done
      -- 
    outputPort_3_Daemon_CP_1538_elements(6) <= outputPort_3_Daemon_CP_1538_elements(158);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	141 
    -- CP-element group 7: 	123 
    -- CP-element group 7: 	21 
    -- CP-element group 7: 	40 
    -- CP-element group 7: 	61 
    -- CP-element group 7: 	82 
    -- CP-element group 7: 	103 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/back_edge_to_loop_body
      -- 
    outputPort_3_Daemon_CP_1538_elements(7) <= outputPort_3_Daemon_CP_1538_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	143 
    -- CP-element group 8: 	125 
    -- CP-element group 8: 	23 
    -- CP-element group 8: 	42 
    -- CP-element group 8: 	63 
    -- CP-element group 8: 	84 
    -- CP-element group 8: 	105 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/first_time_through_loop_body
      -- 
    outputPort_3_Daemon_CP_1538_elements(8) <= outputPort_3_Daemon_CP_1538_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	119 
    -- CP-element group 9: 	157 
    -- CP-element group 9: 	118 
    -- CP-element group 9: 	136 
    -- CP-element group 9: 	137 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	34 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	55 
    -- CP-element group 9: 	56 
    -- CP-element group 9: 	76 
    -- CP-element group 9: 	77 
    -- CP-element group 9: 	97 
    -- CP-element group 9: 	98 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/loop_body_start
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	157 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/condition_evaluated
      -- 
    condition_evaluated_1562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(10), ack => do_while_stmt_1045_branch_req_0); -- 
    outputPort_3_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(157) & outputPort_3_Daemon_CP_1538_elements(14);
      gj_outputPort_3_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	118 
    -- CP-element group 11: 	136 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	55 
    -- CP-element group 11: 	76 
    -- CP-element group 11: 	97 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	138 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	57 
    -- CP-element group 11: 	78 
    -- CP-element group 11: 	99 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1071_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/aggregated_phi_sample_req
      -- 
    outputPort_3_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(118) & outputPort_3_Daemon_CP_1538_elements(136) & outputPort_3_Daemon_CP_1538_elements(15) & outputPort_3_Daemon_CP_1538_elements(34) & outputPort_3_Daemon_CP_1538_elements(55) & outputPort_3_Daemon_CP_1538_elements(76) & outputPort_3_Daemon_CP_1538_elements(97) & outputPort_3_Daemon_CP_1538_elements(14);
      gj_outputPort_3_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	139 
    -- CP-element group 12: 	120 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	37 
    -- CP-element group 12: 	58 
    -- CP-element group 12: 	79 
    -- CP-element group 12: 	100 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	158 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	118 
    -- CP-element group 12: 	136 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	34 
    -- CP-element group 12: 	55 
    -- CP-element group 12: 	76 
    -- CP-element group 12: 	97 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1071_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1075_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1066_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1047_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1051_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1056_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1061_sample_completed_
      -- 
    outputPort_3_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(139) & outputPort_3_Daemon_CP_1538_elements(120) & outputPort_3_Daemon_CP_1538_elements(18) & outputPort_3_Daemon_CP_1538_elements(37) & outputPort_3_Daemon_CP_1538_elements(58) & outputPort_3_Daemon_CP_1538_elements(79) & outputPort_3_Daemon_CP_1538_elements(100);
      gj_outputPort_3_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	119 
    -- CP-element group 13: 	137 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	35 
    -- CP-element group 13: 	56 
    -- CP-element group 13: 	77 
    -- CP-element group 13: 	98 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	121 
    -- CP-element group 13: 	19 
    -- CP-element group 13: 	38 
    -- CP-element group 13: 	59 
    -- CP-element group 13: 	80 
    -- CP-element group 13: 	101 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1075_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/aggregated_phi_update_req
      -- 
    outputPort_3_Daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(119) & outputPort_3_Daemon_CP_1538_elements(137) & outputPort_3_Daemon_CP_1538_elements(16) & outputPort_3_Daemon_CP_1538_elements(35) & outputPort_3_Daemon_CP_1538_elements(56) & outputPort_3_Daemon_CP_1538_elements(77) & outputPort_3_Daemon_CP_1538_elements(98);
      gj_outputPort_3_Daemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	140 
    -- CP-element group 14: 	122 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	60 
    -- CP-element group 14: 	81 
    -- CP-element group 14: 	102 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/aggregated_phi_update_ack
      -- 
    outputPort_3_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(140) & outputPort_3_Daemon_CP_1538_elements(122) & outputPort_3_Daemon_CP_1538_elements(20) & outputPort_3_Daemon_CP_1538_elements(39) & outputPort_3_Daemon_CP_1538_elements(60) & outputPort_3_Daemon_CP_1538_elements(81) & outputPort_3_Daemon_CP_1538_elements(102);
      gj_outputPort_3_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1047_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	155 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1047_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(155);
      gj_outputPort_3_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1047_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(17) <= outputPort_3_Daemon_CP_1538_elements(11);
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1047_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1047_update_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(19) <= outputPort_3_Daemon_CP_1538_elements(13);
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	154 
    -- CP-element group 20: 	14 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1047_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1047_update_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1047_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(21) <= outputPort_3_Daemon_CP_1538_elements(7);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1047_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1047_loopback_sample_req_ps
      -- 
    phi_stmt_1047_loopback_sample_req_1577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1047_loopback_sample_req_1577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(22), ack => phi_stmt_1047_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1047_entry_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(23) <= outputPort_3_Daemon_CP_1538_elements(8);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1047_entry_sample_req
      -- CP-element group 24: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1047_entry_sample_req_ps
      -- 
    phi_stmt_1047_entry_sample_req_1580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1047_entry_sample_req_1580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(24), ack => phi_stmt_1047_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1047_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1047_phi_mux_ack_ps
      -- 
    phi_stmt_1047_phi_mux_ack_1583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1047_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_8_1049_sample_start__ps
      -- CP-element group 26: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_8_1049_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_8_1049_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_8_1049_sample_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_8_1049_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_8_1049_update_start_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_8_1049_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(28) <= outputPort_3_Daemon_CP_1538_elements(29);
    -- CP-element group 29:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	28 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_8_1049_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(29) is a control-delay.
    cp_element_29_delay: control_delay_element  generic map(name => " 29_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_1538_elements(27), ack => outputPort_3_Daemon_CP_1538_elements(29), clk => clk, reset =>reset);
    -- CP-element group 30:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_down_counter_1050_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_down_counter_1050_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_down_counter_1050_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_down_counter_1050_Sample/req
      -- 
    req_1604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(30), ack => next_down_counter_1158_1050_buf_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_down_counter_1050_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_down_counter_1050_update_start_
      -- CP-element group 31: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_down_counter_1050_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_down_counter_1050_Update/req
      -- 
    req_1609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(31), ack => next_down_counter_1158_1050_buf_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_down_counter_1050_sample_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_down_counter_1050_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_down_counter_1050_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_down_counter_1050_Sample/ack
      -- 
    ack_1605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_1158_1050_buf_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(32)); -- 
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_down_counter_1050_update_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_down_counter_1050_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_down_counter_1050_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_down_counter_1050_Update/ack
      -- 
    ack_1610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_1158_1050_buf_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(33)); -- 
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	9 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	12 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	11 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1051_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	155 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	13 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1051_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(155);
      gj_outputPort_3_Daemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	11 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1051_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(36) <= outputPort_3_Daemon_CP_1538_elements(11);
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	12 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1051_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1051_update_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(38) <= outputPort_3_Daemon_CP_1538_elements(13);
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	154 
    -- CP-element group 39: 	14 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1051_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1051_update_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	7 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1051_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(40) <= outputPort_3_Daemon_CP_1538_elements(7);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1051_loopback_sample_req
      -- CP-element group 41: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1051_loopback_sample_req_ps
      -- 
    phi_stmt_1051_loopback_sample_req_1621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1051_loopback_sample_req_1621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(41), ack => phi_stmt_1051_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	8 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1051_entry_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(42) <= outputPort_3_Daemon_CP_1538_elements(8);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1051_entry_sample_req
      -- CP-element group 43: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1051_entry_sample_req_ps
      -- 
    phi_stmt_1051_entry_sample_req_1624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1051_entry_sample_req_1624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(43), ack => phi_stmt_1051_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1051_phi_mux_ack
      -- CP-element group 44: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1051_phi_mux_ack_ps
      -- 
    phi_stmt_1051_phi_mux_ack_1627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1051_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1053_sample_start__ps
      -- CP-element group 45: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1053_sample_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1053_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1053_sample_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1053_update_start__ps
      -- CP-element group 46: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1053_update_start_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1053_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(47) <= outputPort_3_Daemon_CP_1538_elements(48);
    -- CP-element group 48:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	47 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1053_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(48) is a control-delay.
    cp_element_48_delay: control_delay_element  generic map(name => " 48_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_1538_elements(46), ack => outputPort_3_Daemon_CP_1538_elements(48), clk => clk, reset =>reset);
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_1_3_1055_sample_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_1_3_1055_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	54 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_1_3_1055_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_1_3_1055_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_1_3_1055_Sample/rr
      -- 
    rr_1648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(51), ack => RPIPE_noblock_obuf_1_3_1055_inst_req_0); -- 
    outputPort_3_Daemon_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(49) & outputPort_3_Daemon_CP_1538_elements(54);
      gj_outputPort_3_Daemon_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: 	53 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_1_3_1055_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_1_3_1055_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_1_3_1055_Update/cr
      -- 
    cr_1653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(52), ack => RPIPE_noblock_obuf_1_3_1055_inst_req_1); -- 
    outputPort_3_Daemon_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(50) & outputPort_3_Daemon_CP_1538_elements(53);
      gj_outputPort_3_Daemon_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	52 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_1_3_1055_sample_completed__ps
      -- CP-element group 53: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_1_3_1055_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_1_3_1055_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_1_3_1055_Sample/ra
      -- 
    ra_1649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_3_1055_inst_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(53)); -- 
    -- CP-element group 54:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	51 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_1_3_1055_update_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_1_3_1055_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_1_3_1055_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_1_3_1055_Update/ca
      -- 
    ca_1654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_3_1055_inst_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(54)); -- 
    -- CP-element group 55:  join  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	9 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	12 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	11 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1056_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	9 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	155 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	13 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1056_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(155);
      gj_outputPort_3_Daemon_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	11 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1056_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(57) <= outputPort_3_Daemon_CP_1538_elements(11);
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	12 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1056_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	13 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1056_update_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(59) <= outputPort_3_Daemon_CP_1538_elements(13);
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	154 
    -- CP-element group 60: 	14 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1056_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1056_update_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	7 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1056_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(61) <= outputPort_3_Daemon_CP_1538_elements(7);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1056_loopback_sample_req
      -- CP-element group 62: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1056_loopback_sample_req_ps
      -- 
    phi_stmt_1056_loopback_sample_req_1665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1056_loopback_sample_req_1665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(62), ack => phi_stmt_1056_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	8 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1056_entry_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(63) <= outputPort_3_Daemon_CP_1538_elements(8);
    -- CP-element group 64:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1056_entry_sample_req
      -- CP-element group 64: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1056_entry_sample_req_ps
      -- 
    phi_stmt_1056_entry_sample_req_1668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1056_entry_sample_req_1668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(64), ack => phi_stmt_1056_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1056_phi_mux_ack
      -- CP-element group 65: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1056_phi_mux_ack_ps
      -- 
    phi_stmt_1056_phi_mux_ack_1671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1056_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(65)); -- 
    -- CP-element group 66:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1058_sample_start__ps
      -- CP-element group 66: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1058_sample_completed__ps
      -- CP-element group 66: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1058_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1058_sample_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1058_update_start__ps
      -- CP-element group 67: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1058_update_start_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1058_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(68) <= outputPort_3_Daemon_CP_1538_elements(69);
    -- CP-element group 69:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	68 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1058_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(69) is a control-delay.
    cp_element_69_delay: control_delay_element  generic map(name => " 69_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_1538_elements(67), ack => outputPort_3_Daemon_CP_1538_elements(69), clk => clk, reset =>reset);
    -- CP-element group 70:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_2_3_1060_sample_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(70) is bound as output of CP function.
    -- CP-element group 71:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_2_3_1060_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: marked-predecessors 
    -- CP-element group 72: 	75 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_2_3_1060_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_2_3_1060_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_2_3_1060_Sample/rr
      -- 
    rr_1692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(72), ack => RPIPE_noblock_obuf_2_3_1060_inst_req_0); -- 
    outputPort_3_Daemon_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(70) & outputPort_3_Daemon_CP_1538_elements(75);
      gj_outputPort_3_Daemon_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: 	74 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_2_3_1060_update_start_
      -- CP-element group 73: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_2_3_1060_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_2_3_1060_Update/cr
      -- 
    cr_1697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(73), ack => RPIPE_noblock_obuf_2_3_1060_inst_req_1); -- 
    outputPort_3_Daemon_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(71) & outputPort_3_Daemon_CP_1538_elements(74);
      gj_outputPort_3_Daemon_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	73 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_2_3_1060_sample_completed__ps
      -- CP-element group 74: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_2_3_1060_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_2_3_1060_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_2_3_1060_Sample/ra
      -- 
    ra_1693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_3_1060_inst_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(74)); -- 
    -- CP-element group 75:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	72 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_2_3_1060_update_completed__ps
      -- CP-element group 75: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_2_3_1060_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_2_3_1060_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_2_3_1060_Update/ca
      -- 
    ca_1698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_3_1060_inst_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(75)); -- 
    -- CP-element group 76:  join  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	9 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	12 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	11 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1061_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	9 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	155 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	13 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1061_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(155);
      gj_outputPort_3_Daemon_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	11 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1061_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(78) <= outputPort_3_Daemon_CP_1538_elements(11);
    -- CP-element group 79:  join  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	12 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1061_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	13 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1061_update_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(80) <= outputPort_3_Daemon_CP_1538_elements(13);
    -- CP-element group 81:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	154 
    -- CP-element group 81: 	14 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1061_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1061_update_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	7 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1061_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(82) <= outputPort_3_Daemon_CP_1538_elements(7);
    -- CP-element group 83:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1061_loopback_sample_req
      -- CP-element group 83: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1061_loopback_sample_req_ps
      -- 
    phi_stmt_1061_loopback_sample_req_1709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1061_loopback_sample_req_1709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(83), ack => phi_stmt_1061_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(83) is bound as output of CP function.
    -- CP-element group 84:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	8 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1061_entry_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(84) <= outputPort_3_Daemon_CP_1538_elements(8);
    -- CP-element group 85:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1061_entry_sample_req
      -- CP-element group 85: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1061_entry_sample_req_ps
      -- 
    phi_stmt_1061_entry_sample_req_1712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1061_entry_sample_req_1712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(85), ack => phi_stmt_1061_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1061_phi_mux_ack_ps
      -- CP-element group 86: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1061_phi_mux_ack
      -- 
    phi_stmt_1061_phi_mux_ack_1715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1061_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(86)); -- 
    -- CP-element group 87:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1063_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1063_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1063_sample_completed__ps
      -- CP-element group 87: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1063_sample_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1063_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1063_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	90 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1063_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(89) <= outputPort_3_Daemon_CP_1538_elements(90);
    -- CP-element group 90:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	89 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1063_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(90) is a control-delay.
    cp_element_90_delay: control_delay_element  generic map(name => " 90_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_1538_elements(88), ack => outputPort_3_Daemon_CP_1538_elements(90), clk => clk, reset =>reset);
    -- CP-element group 91:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_3_3_1065_sample_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(91) is bound as output of CP function.
    -- CP-element group 92:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_3_3_1065_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(92) is bound as output of CP function.
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	96 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_3_3_1065_Sample/rr
      -- CP-element group 93: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_3_3_1065_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_3_3_1065_sample_start_
      -- 
    rr_1736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(93), ack => RPIPE_noblock_obuf_3_3_1065_inst_req_0); -- 
    outputPort_3_Daemon_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(91) & outputPort_3_Daemon_CP_1538_elements(96);
      gj_outputPort_3_Daemon_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	95 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_3_3_1065_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_3_3_1065_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_3_3_1065_Update/cr
      -- 
    cr_1741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(94), ack => RPIPE_noblock_obuf_3_3_1065_inst_req_1); -- 
    outputPort_3_Daemon_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(92) & outputPort_3_Daemon_CP_1538_elements(95);
      gj_outputPort_3_Daemon_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	94 
    -- CP-element group 95:  members (4) 
      -- CP-element group 95: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_3_3_1065_Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_3_3_1065_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_3_3_1065_sample_completed__ps
      -- CP-element group 95: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_3_3_1065_sample_completed_
      -- 
    ra_1737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_3_1065_inst_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(95)); -- 
    -- CP-element group 96:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	93 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_3_3_1065_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_3_3_1065_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_3_3_1065_Update/ca
      -- CP-element group 96: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_3_3_1065_update_completed__ps
      -- 
    ca_1742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_3_1065_inst_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(96)); -- 
    -- CP-element group 97:  join  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	9 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	12 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	11 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1066_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	9 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	155 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	13 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1066_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(155);
      gj_outputPort_3_Daemon_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	11 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1066_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(99) <= outputPort_3_Daemon_CP_1538_elements(11);
    -- CP-element group 100:  join  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	12 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1066_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(100) is bound as output of CP function.
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	13 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1066_update_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(101) <= outputPort_3_Daemon_CP_1538_elements(13);
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	154 
    -- CP-element group 102: 	14 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1066_update_completed__ps
      -- CP-element group 102: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1066_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(102) is bound as output of CP function.
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	7 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1066_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(103) <= outputPort_3_Daemon_CP_1538_elements(7);
    -- CP-element group 104:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1066_loopback_sample_req_ps
      -- CP-element group 104: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1066_loopback_sample_req
      -- 
    phi_stmt_1066_loopback_sample_req_1753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1066_loopback_sample_req_1753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(104), ack => phi_stmt_1066_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(104) is bound as output of CP function.
    -- CP-element group 105:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	8 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1066_entry_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(105) <= outputPort_3_Daemon_CP_1538_elements(8);
    -- CP-element group 106:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1066_entry_sample_req
      -- CP-element group 106: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1066_entry_sample_req_ps
      -- 
    phi_stmt_1066_entry_sample_req_1756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1066_entry_sample_req_1756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(106), ack => phi_stmt_1066_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1066_phi_mux_ack_ps
      -- CP-element group 107: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1066_phi_mux_ack
      -- 
    phi_stmt_1066_phi_mux_ack_1759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1066_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(107)); -- 
    -- CP-element group 108:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1068_sample_start__ps
      -- CP-element group 108: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1068_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1068_sample_completed__ps
      -- CP-element group 108: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1068_sample_start_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(108) is bound as output of CP function.
    -- CP-element group 109:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1068_update_start__ps
      -- CP-element group 109: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1068_update_start_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	111 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1068_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(110) <= outputPort_3_Daemon_CP_1538_elements(111);
    -- CP-element group 111:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	110 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_33_1068_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(111) is a control-delay.
    cp_element_111_delay: control_delay_element  generic map(name => " 111_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_1538_elements(109), ack => outputPort_3_Daemon_CP_1538_elements(111), clk => clk, reset =>reset);
    -- CP-element group 112:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_4_3_1070_sample_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(112) is bound as output of CP function.
    -- CP-element group 113:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_4_3_1070_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(113) is bound as output of CP function.
    -- CP-element group 114:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: marked-predecessors 
    -- CP-element group 114: 	117 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_4_3_1070_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_4_3_1070_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_4_3_1070_Sample/rr
      -- 
    rr_1780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(114), ack => RPIPE_noblock_obuf_4_3_1070_inst_req_0); -- 
    outputPort_3_Daemon_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(112) & outputPort_3_Daemon_CP_1538_elements(117);
      gj_outputPort_3_Daemon_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	116 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_4_3_1070_Update/cr
      -- CP-element group 115: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_4_3_1070_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_4_3_1070_update_start_
      -- 
    cr_1785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(115), ack => RPIPE_noblock_obuf_4_3_1070_inst_req_1); -- 
    outputPort_3_Daemon_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(113) & outputPort_3_Daemon_CP_1538_elements(116);
      gj_outputPort_3_Daemon_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	115 
    -- CP-element group 116:  members (4) 
      -- CP-element group 116: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_4_3_1070_Sample/ra
      -- CP-element group 116: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_4_3_1070_sample_completed__ps
      -- CP-element group 116: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_4_3_1070_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_4_3_1070_Sample/$exit
      -- 
    ra_1781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_3_1070_inst_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(116)); -- 
    -- CP-element group 117:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: marked-successors 
    -- CP-element group 117: 	114 
    -- CP-element group 117:  members (4) 
      -- CP-element group 117: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_4_3_1070_Update/ca
      -- CP-element group 117: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_4_3_1070_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_4_3_1070_update_completed__ps
      -- CP-element group 117: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/RPIPE_noblock_obuf_4_3_1070_update_completed_
      -- 
    ca_1786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_3_1070_inst_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(117)); -- 
    -- CP-element group 118:  join  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	9 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	12 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	11 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1071_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  join  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	9 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	155 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	13 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1071_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(155);
      gj_outputPort_3_Daemon_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  join  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	12 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1071_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(120) is bound as output of CP function.
    -- CP-element group 121:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	13 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1071_update_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(121) <= outputPort_3_Daemon_CP_1538_elements(13);
    -- CP-element group 122:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	154 
    -- CP-element group 122: 	14 
    -- CP-element group 122:  members (2) 
      -- CP-element group 122: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1071_update_completed__ps
      -- CP-element group 122: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1071_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(122) is bound as output of CP function.
    -- CP-element group 123:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	7 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1071_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(123) <= outputPort_3_Daemon_CP_1538_elements(7);
    -- CP-element group 124:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (2) 
      -- CP-element group 124: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1071_loopback_sample_req
      -- CP-element group 124: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1071_loopback_sample_req_ps
      -- 
    phi_stmt_1071_loopback_sample_req_1797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1071_loopback_sample_req_1797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(124), ack => phi_stmt_1071_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(124) is bound as output of CP function.
    -- CP-element group 125:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	8 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1071_entry_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(125) <= outputPort_3_Daemon_CP_1538_elements(8);
    -- CP-element group 126:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1071_entry_sample_req_ps
      -- CP-element group 126: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1071_entry_sample_req
      -- 
    phi_stmt_1071_entry_sample_req_1800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1071_entry_sample_req_1800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(126), ack => phi_stmt_1071_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(126) is bound as output of CP function.
    -- CP-element group 127:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1071_phi_mux_ack_ps
      -- CP-element group 127: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1071_phi_mux_ack
      -- 
    phi_stmt_1071_phi_mux_ack_1803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1071_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(127)); -- 
    -- CP-element group 128:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (4) 
      -- CP-element group 128: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_3_1073_sample_completed_
      -- CP-element group 128: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_3_1073_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_3_1073_sample_completed__ps
      -- CP-element group 128: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_3_1073_sample_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(128) is bound as output of CP function.
    -- CP-element group 129:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (2) 
      -- CP-element group 129: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_3_1073_update_start_
      -- CP-element group 129: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_3_1073_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(129) is bound as output of CP function.
    -- CP-element group 130:  join  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_3_1073_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(130) <= outputPort_3_Daemon_CP_1538_elements(131);
    -- CP-element group 131:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	130 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ZERO_3_1073_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(131) is a control-delay.
    cp_element_131_delay: control_delay_element  generic map(name => " 131_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_1538_elements(129), ack => outputPort_3_Daemon_CP_1538_elements(131), clk => clk, reset =>reset);
    -- CP-element group 132:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (4) 
      -- CP-element group 132: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_active_packet_1074_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_active_packet_1074_sample_start__ps
      -- CP-element group 132: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_active_packet_1074_Sample/req
      -- CP-element group 132: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_active_packet_1074_sample_start_
      -- 
    req_1824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(132), ack => next_active_packet_1138_1074_buf_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(132) is bound as output of CP function.
    -- CP-element group 133:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	135 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_active_packet_1074_update_start__ps
      -- CP-element group 133: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_active_packet_1074_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_active_packet_1074_Update/req
      -- CP-element group 133: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_active_packet_1074_update_start_
      -- 
    req_1829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(133), ack => next_active_packet_1138_1074_buf_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(133) is bound as output of CP function.
    -- CP-element group 134:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_active_packet_1074_sample_completed__ps
      -- CP-element group 134: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_active_packet_1074_Sample/ack
      -- CP-element group 134: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_active_packet_1074_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_active_packet_1074_Sample/$exit
      -- 
    ack_1825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_1138_1074_buf_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(134)); -- 
    -- CP-element group 135:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	133 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (4) 
      -- CP-element group 135: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_active_packet_1074_Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_active_packet_1074_update_completed__ps
      -- CP-element group 135: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_active_packet_1074_Update/ack
      -- CP-element group 135: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_active_packet_1074_update_completed_
      -- 
    ack_1830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_1138_1074_buf_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(135)); -- 
    -- CP-element group 136:  join  transition  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	9 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	12 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	11 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1075_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  join  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	9 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	155 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	13 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1075_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(155);
      gj_outputPort_3_Daemon_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	11 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1075_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(138) <= outputPort_3_Daemon_CP_1538_elements(11);
    -- CP-element group 139:  join  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	12 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1075_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(139) is bound as output of CP function.
    -- CP-element group 140:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	154 
    -- CP-element group 140: 	14 
    -- CP-element group 140:  members (2) 
      -- CP-element group 140: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1075_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1075_update_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(140) is bound as output of CP function.
    -- CP-element group 141:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	7 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1075_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(141) <= outputPort_3_Daemon_CP_1538_elements(7);
    -- CP-element group 142:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1075_loopback_sample_req
      -- CP-element group 142: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1075_loopback_sample_req_ps
      -- 
    phi_stmt_1075_loopback_sample_req_1841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1075_loopback_sample_req_1841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(142), ack => phi_stmt_1075_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(142) is bound as output of CP function.
    -- CP-element group 143:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	8 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1075_entry_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(143) <= outputPort_3_Daemon_CP_1538_elements(8);
    -- CP-element group 144:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1075_entry_sample_req
      -- CP-element group 144: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1075_entry_sample_req_ps
      -- 
    phi_stmt_1075_entry_sample_req_1844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1075_entry_sample_req_1844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(144), ack => phi_stmt_1075_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1075_phi_mux_ack
      -- CP-element group 145: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/phi_stmt_1075_phi_mux_ack_ps
      -- 
    phi_stmt_1075_phi_mux_ack_1847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1075_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(145)); -- 
    -- CP-element group 146:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (4) 
      -- CP-element group 146: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ONE_3_1077_sample_start__ps
      -- CP-element group 146: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ONE_3_1077_sample_completed__ps
      -- CP-element group 146: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ONE_3_1077_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ONE_3_1077_sample_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(146) is bound as output of CP function.
    -- CP-element group 147:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (2) 
      -- CP-element group 147: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ONE_3_1077_update_start__ps
      -- CP-element group 147: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ONE_3_1077_update_start_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(147) is bound as output of CP function.
    -- CP-element group 148:  join  transition  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	149 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (1) 
      -- CP-element group 148: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ONE_3_1077_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(148) <= outputPort_3_Daemon_CP_1538_elements(149);
    -- CP-element group 149:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	148 
    -- CP-element group 149:  members (1) 
      -- CP-element group 149: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_ONE_3_1077_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(149) is a control-delay.
    cp_element_149_delay: control_delay_element  generic map(name => " 149_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_1538_elements(147), ack => outputPort_3_Daemon_CP_1538_elements(149), clk => clk, reset =>reset);
    -- CP-element group 150:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (4) 
      -- CP-element group 150: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_pkt_priority_1078_Sample/req
      -- CP-element group 150: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_pkt_priority_1078_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_pkt_priority_1078_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_pkt_priority_1078_sample_start__ps
      -- 
    req_1868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(150), ack => next_pkt_priority_1138_1078_buf_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(150) is bound as output of CP function.
    -- CP-element group 151:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (4) 
      -- CP-element group 151: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_pkt_priority_1078_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_pkt_priority_1078_Update/req
      -- CP-element group 151: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_pkt_priority_1078_update_start_
      -- CP-element group 151: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_pkt_priority_1078_update_start__ps
      -- 
    req_1873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(151), ack => next_pkt_priority_1138_1078_buf_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(151) is bound as output of CP function.
    -- CP-element group 152:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (4) 
      -- CP-element group 152: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_pkt_priority_1078_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_pkt_priority_1078_Sample/ack
      -- CP-element group 152: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_pkt_priority_1078_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_pkt_priority_1078_sample_completed__ps
      -- 
    ack_1869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pkt_priority_1138_1078_buf_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(152)); -- 
    -- CP-element group 153:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (4) 
      -- CP-element group 153: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_pkt_priority_1078_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_pkt_priority_1078_Update/ack
      -- CP-element group 153: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_pkt_priority_1078_update_completed__ps
      -- CP-element group 153: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/R_next_pkt_priority_1078_update_completed_
      -- 
    ack_1874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pkt_priority_1138_1078_buf_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	140 
    -- CP-element group 154: 	122 
    -- CP-element group 154: 	20 
    -- CP-element group 154: 	39 
    -- CP-element group 154: 	60 
    -- CP-element group 154: 	81 
    -- CP-element group 154: 	102 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/WPIPE_out_data_3_1265_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/WPIPE_out_data_3_1265_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/WPIPE_out_data_3_1265_Sample/req
      -- 
    req_1883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(154), ack => WPIPE_out_data_3_1265_inst_req_0); -- 
    outputPort_3_Daemon_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(140) & outputPort_3_Daemon_CP_1538_elements(122) & outputPort_3_Daemon_CP_1538_elements(20) & outputPort_3_Daemon_CP_1538_elements(39) & outputPort_3_Daemon_CP_1538_elements(60) & outputPort_3_Daemon_CP_1538_elements(81) & outputPort_3_Daemon_CP_1538_elements(102) & outputPort_3_Daemon_CP_1538_elements(156);
      gj_outputPort_3_Daemon_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	119 
    -- CP-element group 155: 	137 
    -- CP-element group 155: 	16 
    -- CP-element group 155: 	35 
    -- CP-element group 155: 	56 
    -- CP-element group 155: 	77 
    -- CP-element group 155: 	98 
    -- CP-element group 155:  members (6) 
      -- CP-element group 155: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/WPIPE_out_data_3_1265_update_start_
      -- CP-element group 155: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/WPIPE_out_data_3_1265_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/WPIPE_out_data_3_1265_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/WPIPE_out_data_3_1265_Update/req
      -- CP-element group 155: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/WPIPE_out_data_3_1265_Sample/ack
      -- CP-element group 155: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/WPIPE_out_data_3_1265_Update/$entry
      -- 
    ack_1884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_3_1265_inst_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(155)); -- 
    req_1888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(155), ack => WPIPE_out_data_3_1265_inst_req_1); -- 
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	154 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/WPIPE_out_data_3_1265_Update/ack
      -- CP-element group 156: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/WPIPE_out_data_3_1265_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/WPIPE_out_data_3_1265_Update/$exit
      -- 
    ack_1889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_3_1265_inst_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(156)); -- 
    -- CP-element group 157:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	9 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	10 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(157) is a control-delay.
    cp_element_157_delay: control_delay_element  generic map(name => " 157_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_1538_elements(9), ack => outputPort_3_Daemon_CP_1538_elements(157), clk => clk, reset =>reset);
    -- CP-element group 158:  join  transition  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: 	12 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	6 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_1044/do_while_stmt_1045/do_while_stmt_1045_loop_body/$exit
      -- 
    outputPort_3_Daemon_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(156) & outputPort_3_Daemon_CP_1538_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	5 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (2) 
      -- CP-element group 159: 	 branch_block_stmt_1044/do_while_stmt_1045/loop_exit/ack
      -- CP-element group 159: 	 branch_block_stmt_1044/do_while_stmt_1045/loop_exit/$exit
      -- 
    ack_1894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1045_branch_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	5 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (2) 
      -- CP-element group 160: 	 branch_block_stmt_1044/do_while_stmt_1045/loop_taken/$exit
      -- CP-element group 160: 	 branch_block_stmt_1044/do_while_stmt_1045/loop_taken/ack
      -- 
    ack_1898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1045_branch_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(160)); -- 
    -- CP-element group 161:  transition  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	3 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	1 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_1044/do_while_stmt_1045/$exit
      -- 
    outputPort_3_Daemon_CP_1538_elements(161) <= outputPort_3_Daemon_CP_1538_elements(3);
    outputPort_3_Daemon_do_while_stmt_1045_terminator_1899: loop_terminator -- 
      generic map (name => " outputPort_3_Daemon_do_while_stmt_1045_terminator_1899", max_iterations_in_flight =>7) 
      port map(loop_body_exit => outputPort_3_Daemon_CP_1538_elements(6),loop_continue => outputPort_3_Daemon_CP_1538_elements(160),loop_terminate => outputPort_3_Daemon_CP_1538_elements(159),loop_back => outputPort_3_Daemon_CP_1538_elements(4),loop_exit => outputPort_3_Daemon_CP_1538_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1047_phi_seq_1611_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_1538_elements(23);
      outputPort_3_Daemon_CP_1538_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(26);
      outputPort_3_Daemon_CP_1538_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(28);
      outputPort_3_Daemon_CP_1538_elements(24) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_1538_elements(21);
      outputPort_3_Daemon_CP_1538_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(32);
      outputPort_3_Daemon_CP_1538_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(33);
      outputPort_3_Daemon_CP_1538_elements(22) <= phi_mux_reqs(1);
      phi_stmt_1047_phi_seq_1611 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1047_phi_seq_1611") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_1538_elements(17), 
          phi_sample_ack => outputPort_3_Daemon_CP_1538_elements(18), 
          phi_update_req => outputPort_3_Daemon_CP_1538_elements(19), 
          phi_update_ack => outputPort_3_Daemon_CP_1538_elements(20), 
          phi_mux_ack => outputPort_3_Daemon_CP_1538_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1051_phi_seq_1655_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_1538_elements(42);
      outputPort_3_Daemon_CP_1538_elements(45)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(45);
      outputPort_3_Daemon_CP_1538_elements(46)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(47);
      outputPort_3_Daemon_CP_1538_elements(43) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_1538_elements(40);
      outputPort_3_Daemon_CP_1538_elements(49)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(53);
      outputPort_3_Daemon_CP_1538_elements(50)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(54);
      outputPort_3_Daemon_CP_1538_elements(41) <= phi_mux_reqs(1);
      phi_stmt_1051_phi_seq_1655 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1051_phi_seq_1655") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_1538_elements(36), 
          phi_sample_ack => outputPort_3_Daemon_CP_1538_elements(37), 
          phi_update_req => outputPort_3_Daemon_CP_1538_elements(38), 
          phi_update_ack => outputPort_3_Daemon_CP_1538_elements(39), 
          phi_mux_ack => outputPort_3_Daemon_CP_1538_elements(44), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1056_phi_seq_1699_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_1538_elements(63);
      outputPort_3_Daemon_CP_1538_elements(66)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(66);
      outputPort_3_Daemon_CP_1538_elements(67)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(68);
      outputPort_3_Daemon_CP_1538_elements(64) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_1538_elements(61);
      outputPort_3_Daemon_CP_1538_elements(70)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(74);
      outputPort_3_Daemon_CP_1538_elements(71)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(75);
      outputPort_3_Daemon_CP_1538_elements(62) <= phi_mux_reqs(1);
      phi_stmt_1056_phi_seq_1699 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1056_phi_seq_1699") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_1538_elements(57), 
          phi_sample_ack => outputPort_3_Daemon_CP_1538_elements(58), 
          phi_update_req => outputPort_3_Daemon_CP_1538_elements(59), 
          phi_update_ack => outputPort_3_Daemon_CP_1538_elements(60), 
          phi_mux_ack => outputPort_3_Daemon_CP_1538_elements(65), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1061_phi_seq_1743_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_1538_elements(84);
      outputPort_3_Daemon_CP_1538_elements(87)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(87);
      outputPort_3_Daemon_CP_1538_elements(88)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(89);
      outputPort_3_Daemon_CP_1538_elements(85) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_1538_elements(82);
      outputPort_3_Daemon_CP_1538_elements(91)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(95);
      outputPort_3_Daemon_CP_1538_elements(92)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(96);
      outputPort_3_Daemon_CP_1538_elements(83) <= phi_mux_reqs(1);
      phi_stmt_1061_phi_seq_1743 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1061_phi_seq_1743") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_1538_elements(78), 
          phi_sample_ack => outputPort_3_Daemon_CP_1538_elements(79), 
          phi_update_req => outputPort_3_Daemon_CP_1538_elements(80), 
          phi_update_ack => outputPort_3_Daemon_CP_1538_elements(81), 
          phi_mux_ack => outputPort_3_Daemon_CP_1538_elements(86), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1066_phi_seq_1787_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_1538_elements(105);
      outputPort_3_Daemon_CP_1538_elements(108)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(108);
      outputPort_3_Daemon_CP_1538_elements(109)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(110);
      outputPort_3_Daemon_CP_1538_elements(106) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_1538_elements(103);
      outputPort_3_Daemon_CP_1538_elements(112)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(116);
      outputPort_3_Daemon_CP_1538_elements(113)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(117);
      outputPort_3_Daemon_CP_1538_elements(104) <= phi_mux_reqs(1);
      phi_stmt_1066_phi_seq_1787 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1066_phi_seq_1787") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_1538_elements(99), 
          phi_sample_ack => outputPort_3_Daemon_CP_1538_elements(100), 
          phi_update_req => outputPort_3_Daemon_CP_1538_elements(101), 
          phi_update_ack => outputPort_3_Daemon_CP_1538_elements(102), 
          phi_mux_ack => outputPort_3_Daemon_CP_1538_elements(107), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1071_phi_seq_1831_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_1538_elements(125);
      outputPort_3_Daemon_CP_1538_elements(128)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(128);
      outputPort_3_Daemon_CP_1538_elements(129)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(130);
      outputPort_3_Daemon_CP_1538_elements(126) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_1538_elements(123);
      outputPort_3_Daemon_CP_1538_elements(132)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(134);
      outputPort_3_Daemon_CP_1538_elements(133)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(135);
      outputPort_3_Daemon_CP_1538_elements(124) <= phi_mux_reqs(1);
      phi_stmt_1071_phi_seq_1831 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1071_phi_seq_1831") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_1538_elements(11), 
          phi_sample_ack => outputPort_3_Daemon_CP_1538_elements(120), 
          phi_update_req => outputPort_3_Daemon_CP_1538_elements(121), 
          phi_update_ack => outputPort_3_Daemon_CP_1538_elements(122), 
          phi_mux_ack => outputPort_3_Daemon_CP_1538_elements(127), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1075_phi_seq_1875_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_1538_elements(143);
      outputPort_3_Daemon_CP_1538_elements(146)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(146);
      outputPort_3_Daemon_CP_1538_elements(147)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(148);
      outputPort_3_Daemon_CP_1538_elements(144) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_1538_elements(141);
      outputPort_3_Daemon_CP_1538_elements(150)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(152);
      outputPort_3_Daemon_CP_1538_elements(151)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(153);
      outputPort_3_Daemon_CP_1538_elements(142) <= phi_mux_reqs(1);
      phi_stmt_1075_phi_seq_1875 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1075_phi_seq_1875") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_1538_elements(138), 
          phi_sample_ack => outputPort_3_Daemon_CP_1538_elements(139), 
          phi_update_req => outputPort_3_Daemon_CP_1538_elements(13), 
          phi_update_ack => outputPort_3_Daemon_CP_1538_elements(140), 
          phi_mux_ack => outputPort_3_Daemon_CP_1538_elements(145), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1563_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= outputPort_3_Daemon_CP_1538_elements(7);
        preds(1)  <= outputPort_3_Daemon_CP_1538_elements(8);
        entry_tmerge_1563 : transition_merge -- 
          generic map(name => " entry_tmerge_1563")
          port map (preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u3_u1_1103_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1109_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1116_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1122_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1164_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1172_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1180_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1188_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1205_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1212_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1220_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1227_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1238_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1244_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1251_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1257_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_1145_wire : std_logic_vector(0 downto 0);
    signal MUX_1106_wire : std_logic_vector(0 downto 0);
    signal MUX_1112_wire : std_logic_vector(0 downto 0);
    signal MUX_1119_wire : std_logic_vector(0 downto 0);
    signal MUX_1125_wire : std_logic_vector(0 downto 0);
    signal MUX_1156_wire : std_logic_vector(7 downto 0);
    signal MUX_1209_wire : std_logic_vector(31 downto 0);
    signal MUX_1216_wire : std_logic_vector(31 downto 0);
    signal MUX_1224_wire : std_logic_vector(31 downto 0);
    signal MUX_1231_wire : std_logic_vector(31 downto 0);
    signal MUX_1241_wire : std_logic_vector(0 downto 0);
    signal MUX_1247_wire : std_logic_vector(0 downto 0);
    signal MUX_1254_wire : std_logic_vector(0 downto 0);
    signal MUX_1260_wire : std_logic_vector(0 downto 0);
    signal NEQ_u3_u1_1142_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1161_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1169_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1177_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1185_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1113_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1126_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1248_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1261_wire : std_logic_vector(0 downto 0);
    signal OR_u32_u32_1217_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_1232_wire : std_logic_vector(31 downto 0);
    signal RPIPE_noblock_obuf_1_3_1055_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_2_3_1060_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_3_3_1065_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_4_3_1070_wire : std_logic_vector(32 downto 0);
    signal R_ONE_3_1077_wire_constant : std_logic_vector(2 downto 0);
    signal R_ZERO_33_1053_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1058_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1063_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1068_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_3_1073_wire_constant : std_logic_vector(2 downto 0);
    signal R_ZERO_8_1049_wire_constant : std_logic_vector(7 downto 0);
    signal SUB_u8_u8_1154_wire : std_logic_vector(7 downto 0);
    signal active_packet_1071 : std_logic_vector(2 downto 0);
    signal data_to_out_1234 : std_logic_vector(31 downto 0);
    signal down_counter_1047 : std_logic_vector(7 downto 0);
    signal konst_1082_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1087_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1092_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1097_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1102_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1105_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1108_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1111_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1115_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1118_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1121_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1124_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1141_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1144_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1150_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1153_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1163_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1171_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1179_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1187_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1204_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1208_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1211_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1215_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1219_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1223_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1226_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1230_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1237_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1240_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1243_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1246_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1250_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1253_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1256_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1259_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1269_wire_constant : std_logic_vector(0 downto 0);
    signal next_active_packet_1138 : std_logic_vector(2 downto 0);
    signal next_active_packet_1138_1074_buffered : std_logic_vector(2 downto 0);
    signal next_down_counter_1158 : std_logic_vector(7 downto 0);
    signal next_down_counter_1158_1050_buffered : std_logic_vector(7 downto 0);
    signal next_pkt_priority_1138 : std_logic_vector(2 downto 0);
    signal next_pkt_priority_1138_1078_buffered : std_logic_vector(2 downto 0);
    signal p1_valid_1084 : std_logic_vector(0 downto 0);
    signal p2_valid_1089 : std_logic_vector(0 downto 0);
    signal p3_valid_1094 : std_logic_vector(0 downto 0);
    signal p4_valid_1099 : std_logic_vector(0 downto 0);
    signal pkt_1_e_word_1051 : std_logic_vector(32 downto 0);
    signal pkt_2_e_word_1056 : std_logic_vector(32 downto 0);
    signal pkt_3_e_word_1061 : std_logic_vector(32 downto 0);
    signal pkt_4_e_word_1066 : std_logic_vector(32 downto 0);
    signal pkt_priority_1075 : std_logic_vector(2 downto 0);
    signal read_from_1_1166 : std_logic_vector(0 downto 0);
    signal read_from_2_1174 : std_logic_vector(0 downto 0);
    signal read_from_3_1182 : std_logic_vector(0 downto 0);
    signal read_from_4_1190 : std_logic_vector(0 downto 0);
    signal send_flag_1263 : std_logic_vector(0 downto 0);
    signal slice_1207_wire : std_logic_vector(31 downto 0);
    signal slice_1214_wire : std_logic_vector(31 downto 0);
    signal slice_1222_wire : std_logic_vector(31 downto 0);
    signal slice_1229_wire : std_logic_vector(31 downto 0);
    signal started_new_packet_1147 : std_logic_vector(0 downto 0);
    signal valid_active_pkt_word_read_1128 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_ONE_3_1077_wire_constant <= "001";
    R_ZERO_33_1053_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1058_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1063_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1068_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_3_1073_wire_constant <= "000";
    R_ZERO_8_1049_wire_constant <= "00000000";
    konst_1082_wire_constant <= "000000000000000000000000000100000";
    konst_1087_wire_constant <= "000000000000000000000000000100000";
    konst_1092_wire_constant <= "000000000000000000000000000100000";
    konst_1097_wire_constant <= "000000000000000000000000000100000";
    konst_1102_wire_constant <= "001";
    konst_1105_wire_constant <= "0";
    konst_1108_wire_constant <= "010";
    konst_1111_wire_constant <= "0";
    konst_1115_wire_constant <= "011";
    konst_1118_wire_constant <= "0";
    konst_1121_wire_constant <= "100";
    konst_1124_wire_constant <= "0";
    konst_1141_wire_constant <= "000";
    konst_1144_wire_constant <= "00000000";
    konst_1150_wire_constant <= "00111111";
    konst_1153_wire_constant <= "00000001";
    konst_1163_wire_constant <= "001";
    konst_1171_wire_constant <= "010";
    konst_1179_wire_constant <= "011";
    konst_1187_wire_constant <= "100";
    konst_1204_wire_constant <= "001";
    konst_1208_wire_constant <= "00000000000000000000000000000000";
    konst_1211_wire_constant <= "010";
    konst_1215_wire_constant <= "00000000000000000000000000000000";
    konst_1219_wire_constant <= "011";
    konst_1223_wire_constant <= "00000000000000000000000000000000";
    konst_1226_wire_constant <= "100";
    konst_1230_wire_constant <= "00000000000000000000000000000000";
    konst_1237_wire_constant <= "001";
    konst_1240_wire_constant <= "0";
    konst_1243_wire_constant <= "010";
    konst_1246_wire_constant <= "0";
    konst_1250_wire_constant <= "011";
    konst_1253_wire_constant <= "0";
    konst_1256_wire_constant <= "100";
    konst_1259_wire_constant <= "0";
    konst_1269_wire_constant <= "1";
    phi_stmt_1047: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_8_1049_wire_constant & next_down_counter_1158_1050_buffered;
      req <= phi_stmt_1047_req_0 & phi_stmt_1047_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1047",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1047_ack_0,
          idata => idata,
          odata => down_counter_1047,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1047
    phi_stmt_1051: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1053_wire_constant & RPIPE_noblock_obuf_1_3_1055_wire;
      req <= phi_stmt_1051_req_0 & phi_stmt_1051_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1051",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1051_ack_0,
          idata => idata,
          odata => pkt_1_e_word_1051,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1051
    phi_stmt_1056: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1058_wire_constant & RPIPE_noblock_obuf_2_3_1060_wire;
      req <= phi_stmt_1056_req_0 & phi_stmt_1056_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1056",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1056_ack_0,
          idata => idata,
          odata => pkt_2_e_word_1056,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1056
    phi_stmt_1061: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1063_wire_constant & RPIPE_noblock_obuf_3_3_1065_wire;
      req <= phi_stmt_1061_req_0 & phi_stmt_1061_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1061",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1061_ack_0,
          idata => idata,
          odata => pkt_3_e_word_1061,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1061
    phi_stmt_1066: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1068_wire_constant & RPIPE_noblock_obuf_4_3_1070_wire;
      req <= phi_stmt_1066_req_0 & phi_stmt_1066_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1066",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1066_ack_0,
          idata => idata,
          odata => pkt_4_e_word_1066,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1066
    phi_stmt_1071: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_3_1073_wire_constant & next_active_packet_1138_1074_buffered;
      req <= phi_stmt_1071_req_0 & phi_stmt_1071_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1071",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1071_ack_0,
          idata => idata,
          odata => active_packet_1071,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1071
    phi_stmt_1075: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ONE_3_1077_wire_constant & next_pkt_priority_1138_1078_buffered;
      req <= phi_stmt_1075_req_0 & phi_stmt_1075_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1075",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1075_ack_0,
          idata => idata,
          odata => pkt_priority_1075,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1075
    -- flow-through select operator MUX_1106_inst
    MUX_1106_wire <= p1_valid_1084 when (EQ_u3_u1_1103_wire(0) /=  '0') else konst_1105_wire_constant;
    -- flow-through select operator MUX_1112_inst
    MUX_1112_wire <= p2_valid_1089 when (EQ_u3_u1_1109_wire(0) /=  '0') else konst_1111_wire_constant;
    -- flow-through select operator MUX_1119_inst
    MUX_1119_wire <= p3_valid_1094 when (EQ_u3_u1_1116_wire(0) /=  '0') else konst_1118_wire_constant;
    -- flow-through select operator MUX_1125_inst
    MUX_1125_wire <= p4_valid_1099 when (EQ_u3_u1_1122_wire(0) /=  '0') else konst_1124_wire_constant;
    -- flow-through select operator MUX_1156_inst
    MUX_1156_wire <= SUB_u8_u8_1154_wire when (valid_active_pkt_word_read_1128(0) /=  '0') else down_counter_1047;
    -- flow-through select operator MUX_1157_inst
    next_down_counter_1158 <= konst_1150_wire_constant when (started_new_packet_1147(0) /=  '0') else MUX_1156_wire;
    -- flow-through select operator MUX_1209_inst
    MUX_1209_wire <= slice_1207_wire when (EQ_u3_u1_1205_wire(0) /=  '0') else konst_1208_wire_constant;
    -- flow-through select operator MUX_1216_inst
    MUX_1216_wire <= slice_1214_wire when (EQ_u3_u1_1212_wire(0) /=  '0') else konst_1215_wire_constant;
    -- flow-through select operator MUX_1224_inst
    MUX_1224_wire <= slice_1222_wire when (EQ_u3_u1_1220_wire(0) /=  '0') else konst_1223_wire_constant;
    -- flow-through select operator MUX_1231_inst
    MUX_1231_wire <= slice_1229_wire when (EQ_u3_u1_1227_wire(0) /=  '0') else konst_1230_wire_constant;
    -- flow-through select operator MUX_1241_inst
    MUX_1241_wire <= p1_valid_1084 when (EQ_u3_u1_1238_wire(0) /=  '0') else konst_1240_wire_constant;
    -- flow-through select operator MUX_1247_inst
    MUX_1247_wire <= p2_valid_1089 when (EQ_u3_u1_1244_wire(0) /=  '0') else konst_1246_wire_constant;
    -- flow-through select operator MUX_1254_inst
    MUX_1254_wire <= p3_valid_1094 when (EQ_u3_u1_1251_wire(0) /=  '0') else konst_1253_wire_constant;
    -- flow-through select operator MUX_1260_inst
    MUX_1260_wire <= p4_valid_1099 when (EQ_u3_u1_1257_wire(0) /=  '0') else konst_1259_wire_constant;
    -- flow-through slice operator slice_1207_inst
    slice_1207_wire <= pkt_1_e_word_1051(31 downto 0);
    -- flow-through slice operator slice_1214_inst
    slice_1214_wire <= pkt_2_e_word_1056(31 downto 0);
    -- flow-through slice operator slice_1222_inst
    slice_1222_wire <= pkt_3_e_word_1061(31 downto 0);
    -- flow-through slice operator slice_1229_inst
    slice_1229_wire <= pkt_4_e_word_1066(31 downto 0);
    next_active_packet_1138_1074_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_active_packet_1138_1074_buf_req_0;
      next_active_packet_1138_1074_buf_ack_0<= wack(0);
      rreq(0) <= next_active_packet_1138_1074_buf_req_1;
      next_active_packet_1138_1074_buf_ack_1<= rack(0);
      next_active_packet_1138_1074_buf : InterlockBuffer generic map ( -- 
        name => "next_active_packet_1138_1074_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_active_packet_1138,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_active_packet_1138_1074_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_down_counter_1158_1050_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_down_counter_1158_1050_buf_req_0;
      next_down_counter_1158_1050_buf_ack_0<= wack(0);
      rreq(0) <= next_down_counter_1158_1050_buf_req_1;
      next_down_counter_1158_1050_buf_ack_1<= rack(0);
      next_down_counter_1158_1050_buf : InterlockBuffer generic map ( -- 
        name => "next_down_counter_1158_1050_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_down_counter_1158,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_down_counter_1158_1050_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_pkt_priority_1138_1078_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_pkt_priority_1138_1078_buf_req_0;
      next_pkt_priority_1138_1078_buf_ack_0<= wack(0);
      rreq(0) <= next_pkt_priority_1138_1078_buf_req_1;
      next_pkt_priority_1138_1078_buf_ack_1<= rack(0);
      next_pkt_priority_1138_1078_buf : InterlockBuffer generic map ( -- 
        name => "next_pkt_priority_1138_1078_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_pkt_priority_1138,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_pkt_priority_1138_1078_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1045_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1269_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1045_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1045_branch_req_0,
          ack0 => do_while_stmt_1045_branch_ack_0,
          ack1 => do_while_stmt_1045_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator AND_u1_u1_1146_inst
    process(NEQ_u3_u1_1142_wire, EQ_u8_u1_1145_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NEQ_u3_u1_1142_wire, EQ_u8_u1_1145_wire, tmp_var);
      started_new_packet_1147 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_1083_inst
    process(pkt_1_e_word_1051) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_1_e_word_1051, konst_1082_wire_constant, tmp_var);
      p1_valid_1084 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_1088_inst
    process(pkt_2_e_word_1056) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_2_e_word_1056, konst_1087_wire_constant, tmp_var);
      p2_valid_1089 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_1093_inst
    process(pkt_3_e_word_1061) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_3_e_word_1061, konst_1092_wire_constant, tmp_var);
      p3_valid_1094 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_1098_inst
    process(pkt_4_e_word_1066) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_4_e_word_1066, konst_1097_wire_constant, tmp_var);
      p4_valid_1099 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1103_inst
    process(active_packet_1071) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1071, konst_1102_wire_constant, tmp_var);
      EQ_u3_u1_1103_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1109_inst
    process(active_packet_1071) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1071, konst_1108_wire_constant, tmp_var);
      EQ_u3_u1_1109_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1116_inst
    process(active_packet_1071) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1071, konst_1115_wire_constant, tmp_var);
      EQ_u3_u1_1116_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1122_inst
    process(active_packet_1071) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1071, konst_1121_wire_constant, tmp_var);
      EQ_u3_u1_1122_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1164_inst
    process(next_active_packet_1138) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1138, konst_1163_wire_constant, tmp_var);
      EQ_u3_u1_1164_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1172_inst
    process(next_active_packet_1138) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1138, konst_1171_wire_constant, tmp_var);
      EQ_u3_u1_1172_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1180_inst
    process(next_active_packet_1138) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1138, konst_1179_wire_constant, tmp_var);
      EQ_u3_u1_1180_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1188_inst
    process(next_active_packet_1138) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1138, konst_1187_wire_constant, tmp_var);
      EQ_u3_u1_1188_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1205_inst
    process(next_active_packet_1138) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1138, konst_1204_wire_constant, tmp_var);
      EQ_u3_u1_1205_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1212_inst
    process(next_active_packet_1138) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1138, konst_1211_wire_constant, tmp_var);
      EQ_u3_u1_1212_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1220_inst
    process(next_active_packet_1138) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1138, konst_1219_wire_constant, tmp_var);
      EQ_u3_u1_1220_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1227_inst
    process(next_active_packet_1138) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1138, konst_1226_wire_constant, tmp_var);
      EQ_u3_u1_1227_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1238_inst
    process(next_active_packet_1138) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1138, konst_1237_wire_constant, tmp_var);
      EQ_u3_u1_1238_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1244_inst
    process(next_active_packet_1138) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1138, konst_1243_wire_constant, tmp_var);
      EQ_u3_u1_1244_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1251_inst
    process(next_active_packet_1138) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1138, konst_1250_wire_constant, tmp_var);
      EQ_u3_u1_1251_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1257_inst
    process(next_active_packet_1138) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1138, konst_1256_wire_constant, tmp_var);
      EQ_u3_u1_1257_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_1145_inst
    process(down_counter_1047) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(down_counter_1047, konst_1144_wire_constant, tmp_var);
      EQ_u8_u1_1145_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u3_u1_1142_inst
    process(next_active_packet_1138) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(next_active_packet_1138, konst_1141_wire_constant, tmp_var);
      NEQ_u3_u1_1142_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1161_inst
    process(p1_valid_1084) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_1084, tmp_var);
      NOT_u1_u1_1161_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1169_inst
    process(p2_valid_1089) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_1089, tmp_var);
      NOT_u1_u1_1169_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1177_inst
    process(p3_valid_1094) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_1094, tmp_var);
      NOT_u1_u1_1177_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1185_inst
    process(p4_valid_1099) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_1099, tmp_var);
      NOT_u1_u1_1185_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1113_inst
    process(MUX_1106_wire, MUX_1112_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1106_wire, MUX_1112_wire, tmp_var);
      OR_u1_u1_1113_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1126_inst
    process(MUX_1119_wire, MUX_1125_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1119_wire, MUX_1125_wire, tmp_var);
      OR_u1_u1_1126_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1127_inst
    process(OR_u1_u1_1113_wire, OR_u1_u1_1126_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1113_wire, OR_u1_u1_1126_wire, tmp_var);
      valid_active_pkt_word_read_1128 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1165_inst
    process(NOT_u1_u1_1161_wire, EQ_u3_u1_1164_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1161_wire, EQ_u3_u1_1164_wire, tmp_var);
      read_from_1_1166 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1173_inst
    process(NOT_u1_u1_1169_wire, EQ_u3_u1_1172_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1169_wire, EQ_u3_u1_1172_wire, tmp_var);
      read_from_2_1174 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1181_inst
    process(NOT_u1_u1_1177_wire, EQ_u3_u1_1180_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1177_wire, EQ_u3_u1_1180_wire, tmp_var);
      read_from_3_1182 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1189_inst
    process(NOT_u1_u1_1185_wire, EQ_u3_u1_1188_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1185_wire, EQ_u3_u1_1188_wire, tmp_var);
      read_from_4_1190 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1248_inst
    process(MUX_1241_wire, MUX_1247_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1241_wire, MUX_1247_wire, tmp_var);
      OR_u1_u1_1248_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1261_inst
    process(MUX_1254_wire, MUX_1260_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1254_wire, MUX_1260_wire, tmp_var);
      OR_u1_u1_1261_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1262_inst
    process(OR_u1_u1_1248_wire, OR_u1_u1_1261_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1248_wire, OR_u1_u1_1261_wire, tmp_var);
      send_flag_1263 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1217_inst
    process(MUX_1209_wire, MUX_1216_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1209_wire, MUX_1216_wire, tmp_var);
      OR_u32_u32_1217_wire <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1232_inst
    process(MUX_1224_wire, MUX_1231_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1224_wire, MUX_1231_wire, tmp_var);
      OR_u32_u32_1232_wire <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1233_inst
    process(OR_u32_u32_1217_wire, OR_u32_u32_1232_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u32_u32_1217_wire, OR_u32_u32_1232_wire, tmp_var);
      data_to_out_1234 <= tmp_var; --
    end process;
    -- binary operator SUB_u8_u8_1154_inst
    process(down_counter_1047) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSub_proc(down_counter_1047, konst_1153_wire_constant, tmp_var);
      SUB_u8_u8_1154_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_noblock_obuf_1_3_1055_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_1_3_1055_inst_req_0;
      RPIPE_noblock_obuf_1_3_1055_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_1_3_1055_inst_req_1;
      RPIPE_noblock_obuf_1_3_1055_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_1_1166(0);
      RPIPE_noblock_obuf_1_3_1055_wire <= data_out(32 downto 0);
      noblock_obuf_1_3_read_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_3_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_3_read_0: InputPortRevised -- 
        generic map ( name => "noblock_obuf_1_3_read_0", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_1_3_pipe_read_req(0),
          oack => noblock_obuf_1_3_pipe_read_ack(0),
          odata => noblock_obuf_1_3_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_noblock_obuf_2_3_1060_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_2_3_1060_inst_req_0;
      RPIPE_noblock_obuf_2_3_1060_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_2_3_1060_inst_req_1;
      RPIPE_noblock_obuf_2_3_1060_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_2_1174(0);
      RPIPE_noblock_obuf_2_3_1060_wire <= data_out(32 downto 0);
      noblock_obuf_2_3_read_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_3_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_3_read_1: InputPortRevised -- 
        generic map ( name => "noblock_obuf_2_3_read_1", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_2_3_pipe_read_req(0),
          oack => noblock_obuf_2_3_pipe_read_ack(0),
          odata => noblock_obuf_2_3_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_noblock_obuf_3_3_1065_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_3_3_1065_inst_req_0;
      RPIPE_noblock_obuf_3_3_1065_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_3_3_1065_inst_req_1;
      RPIPE_noblock_obuf_3_3_1065_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_3_1182(0);
      RPIPE_noblock_obuf_3_3_1065_wire <= data_out(32 downto 0);
      noblock_obuf_3_3_read_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_3_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_3_read_2: InputPortRevised -- 
        generic map ( name => "noblock_obuf_3_3_read_2", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_3_3_pipe_read_req(0),
          oack => noblock_obuf_3_3_pipe_read_ack(0),
          odata => noblock_obuf_3_3_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_noblock_obuf_4_3_1070_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_4_3_1070_inst_req_0;
      RPIPE_noblock_obuf_4_3_1070_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_4_3_1070_inst_req_1;
      RPIPE_noblock_obuf_4_3_1070_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_4_1190(0);
      RPIPE_noblock_obuf_4_3_1070_wire <= data_out(32 downto 0);
      noblock_obuf_4_3_read_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_3_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_3_read_3: InputPortRevised -- 
        generic map ( name => "noblock_obuf_4_3_read_3", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_4_3_pipe_read_req(0),
          oack => noblock_obuf_4_3_pipe_read_ack(0),
          odata => noblock_obuf_4_3_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_out_data_3_1265_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_out_data_3_1265_inst_req_0;
      WPIPE_out_data_3_1265_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_out_data_3_1265_inst_req_1;
      WPIPE_out_data_3_1265_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_flag_1263(0);
      data_in <= data_to_out_1234;
      out_data_3_write_0_gI: SplitGuardInterface generic map(name => "out_data_3_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      out_data_3_write_0: OutputPortRevised -- 
        generic map ( name => "out_data_3", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => out_data_3_pipe_write_req(0),
          oack => out_data_3_pipe_write_ack(0),
          odata => out_data_3_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    volatile_operator_prioritySelect_3080: prioritySelect_Volatile port map(down_counter => down_counter_1047, active_packet => active_packet_1071, pkt_priority => pkt_priority_1075, p1_valid => p1_valid_1084, p2_valid => p2_valid_1089, p3_valid => p3_valid_1094, p4_valid => p4_valid_1099, next_active_packet => next_active_packet_1138, next_pkt_priority => next_pkt_priority_1138); 
    -- 
  end Block; -- data_path
  -- 
end outputPort_3_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity outputPort_4_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    noblock_obuf_1_4_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_4_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_3_4_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_4_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_2_4_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_4_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_4_4_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_4_pipe_read_data : in   std_logic_vector(32 downto 0);
    out_data_4_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_4_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity outputPort_4_Daemon;
architecture outputPort_4_Daemon_arch of outputPort_4_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal outputPort_4_Daemon_CP_1900_start: Boolean;
  signal outputPort_4_Daemon_CP_1900_symbol: Boolean;
  -- volatile/operator module components. 
  component prioritySelect_Volatile is -- 
    port ( -- 
      down_counter : in  std_logic_vector(7 downto 0);
      active_packet : in  std_logic_vector(2 downto 0);
      pkt_priority : in  std_logic_vector(2 downto 0);
      p1_valid : in  std_logic_vector(0 downto 0);
      p2_valid : in  std_logic_vector(0 downto 0);
      p3_valid : in  std_logic_vector(0 downto 0);
      p4_valid : in  std_logic_vector(0 downto 0);
      next_active_packet : out  std_logic_vector(2 downto 0);
      next_pkt_priority : out  std_logic_vector(2 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal RPIPE_noblock_obuf_3_4_1294_inst_ack_1 : boolean;
  signal RPIPE_noblock_obuf_3_4_1294_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_3_4_1294_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_1_4_1284_inst_ack_1 : boolean;
  signal RPIPE_noblock_obuf_3_4_1294_inst_ack_0 : boolean;
  signal phi_stmt_1290_req_0 : boolean;
  signal phi_stmt_1300_ack_0 : boolean;
  signal phi_stmt_1295_req_0 : boolean;
  signal WPIPE_out_data_4_1494_inst_req_1 : boolean;
  signal next_pkt_priority_1367_1307_buf_ack_1 : boolean;
  signal next_active_packet_1367_1303_buf_req_0 : boolean;
  signal next_pkt_priority_1367_1307_buf_req_1 : boolean;
  signal phi_stmt_1300_req_0 : boolean;
  signal phi_stmt_1290_req_1 : boolean;
  signal RPIPE_noblock_obuf_1_4_1284_inst_req_0 : boolean;
  signal next_active_packet_1367_1303_buf_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_4_1284_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_4_1284_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_2_4_1289_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_2_4_1289_inst_ack_0 : boolean;
  signal phi_stmt_1300_req_1 : boolean;
  signal RPIPE_noblock_obuf_2_4_1289_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_2_4_1289_inst_ack_1 : boolean;
  signal RPIPE_noblock_obuf_4_4_1299_inst_req_1 : boolean;
  signal phi_stmt_1295_req_1 : boolean;
  signal phi_stmt_1295_ack_0 : boolean;
  signal RPIPE_noblock_obuf_4_4_1299_inst_req_0 : boolean;
  signal next_pkt_priority_1367_1307_buf_ack_0 : boolean;
  signal next_pkt_priority_1367_1307_buf_req_0 : boolean;
  signal WPIPE_out_data_4_1494_inst_ack_0 : boolean;
  signal WPIPE_out_data_4_1494_inst_req_0 : boolean;
  signal WPIPE_out_data_4_1494_inst_ack_1 : boolean;
  signal phi_stmt_1280_ack_0 : boolean;
  signal RPIPE_noblock_obuf_4_4_1299_inst_ack_1 : boolean;
  signal phi_stmt_1285_ack_0 : boolean;
  signal phi_stmt_1285_req_0 : boolean;
  signal next_active_packet_1367_1303_buf_ack_1 : boolean;
  signal phi_stmt_1285_req_1 : boolean;
  signal next_active_packet_1367_1303_buf_req_1 : boolean;
  signal phi_stmt_1304_ack_0 : boolean;
  signal phi_stmt_1290_ack_0 : boolean;
  signal phi_stmt_1304_req_0 : boolean;
  signal phi_stmt_1304_req_1 : boolean;
  signal do_while_stmt_1274_branch_req_0 : boolean;
  signal phi_stmt_1276_req_1 : boolean;
  signal phi_stmt_1276_req_0 : boolean;
  signal phi_stmt_1276_ack_0 : boolean;
  signal RPIPE_noblock_obuf_4_4_1299_inst_ack_0 : boolean;
  signal next_down_counter_1387_1279_buf_req_0 : boolean;
  signal next_down_counter_1387_1279_buf_ack_0 : boolean;
  signal next_down_counter_1387_1279_buf_req_1 : boolean;
  signal next_down_counter_1387_1279_buf_ack_1 : boolean;
  signal phi_stmt_1280_req_1 : boolean;
  signal phi_stmt_1280_req_0 : boolean;
  signal do_while_stmt_1274_branch_ack_0 : boolean;
  signal do_while_stmt_1274_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "outputPort_4_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  outputPort_4_Daemon_CP_1900_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "outputPort_4_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_4_Daemon_CP_1900_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= outputPort_4_Daemon_CP_1900_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_4_Daemon_CP_1900_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  outputPort_4_Daemon_CP_1900: Block -- control-path 
    signal outputPort_4_Daemon_CP_1900_elements: BooleanArray(161 downto 0);
    -- 
  begin -- 
    outputPort_4_Daemon_CP_1900_elements(0) <= outputPort_4_Daemon_CP_1900_start;
    outputPort_4_Daemon_CP_1900_symbol <= outputPort_4_Daemon_CP_1900_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1273/$entry
      -- CP-element group 0: 	 branch_block_stmt_1273/branch_block_stmt_1273__entry__
      -- CP-element group 0: 	 branch_block_stmt_1273/do_while_stmt_1274__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	161 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1273/$exit
      -- CP-element group 1: 	 branch_block_stmt_1273/branch_block_stmt_1273__exit__
      -- CP-element group 1: 	 branch_block_stmt_1273/do_while_stmt_1274__exit__
      -- 
    outputPort_4_Daemon_CP_1900_elements(1) <= outputPort_4_Daemon_CP_1900_elements(161);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1273/do_while_stmt_1274/$entry
      -- CP-element group 2: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274__entry__
      -- 
    outputPort_4_Daemon_CP_1900_elements(2) <= outputPort_4_Daemon_CP_1900_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	161 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274__exit__
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1273/do_while_stmt_1274/loop_back
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	159 
    -- CP-element group 5: 	160 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1273/do_while_stmt_1274/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1273/do_while_stmt_1274/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1273/do_while_stmt_1274/loop_taken/$entry
      -- 
    outputPort_4_Daemon_CP_1900_elements(5) <= outputPort_4_Daemon_CP_1900_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	158 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1273/do_while_stmt_1274/loop_body_done
      -- 
    outputPort_4_Daemon_CP_1900_elements(6) <= outputPort_4_Daemon_CP_1900_elements(158);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	141 
    -- CP-element group 7: 	82 
    -- CP-element group 7: 	123 
    -- CP-element group 7: 	102 
    -- CP-element group 7: 	21 
    -- CP-element group 7: 	40 
    -- CP-element group 7: 	61 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/back_edge_to_loop_body
      -- 
    outputPort_4_Daemon_CP_1900_elements(7) <= outputPort_4_Daemon_CP_1900_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	125 
    -- CP-element group 8: 	104 
    -- CP-element group 8: 	143 
    -- CP-element group 8: 	84 
    -- CP-element group 8: 	23 
    -- CP-element group 8: 	42 
    -- CP-element group 8: 	63 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/first_time_through_loop_body
      -- 
    outputPort_4_Daemon_CP_1900_elements(8) <= outputPort_4_Daemon_CP_1900_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	98 
    -- CP-element group 9: 	117 
    -- CP-element group 9: 	136 
    -- CP-element group 9: 	137 
    -- CP-element group 9: 	97 
    -- CP-element group 9: 	118 
    -- CP-element group 9: 	157 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	34 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	55 
    -- CP-element group 9: 	56 
    -- CP-element group 9: 	76 
    -- CP-element group 9: 	77 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/loop_body_start
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	157 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/condition_evaluated
      -- 
    condition_evaluated_1924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(10), ack => do_while_stmt_1274_branch_req_0); -- 
    outputPort_4_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(157) & outputPort_4_Daemon_CP_1900_elements(14);
      gj_outputPort_4_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	117 
    -- CP-element group 11: 	136 
    -- CP-element group 11: 	97 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	55 
    -- CP-element group 11: 	76 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	138 
    -- CP-element group 11: 	119 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	57 
    -- CP-element group 11: 	78 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1295_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/aggregated_phi_sample_req
      -- 
    outputPort_4_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(117) & outputPort_4_Daemon_CP_1900_elements(136) & outputPort_4_Daemon_CP_1900_elements(97) & outputPort_4_Daemon_CP_1900_elements(15) & outputPort_4_Daemon_CP_1900_elements(34) & outputPort_4_Daemon_CP_1900_elements(55) & outputPort_4_Daemon_CP_1900_elements(76) & outputPort_4_Daemon_CP_1900_elements(14);
      gj_outputPort_4_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	139 
    -- CP-element group 12: 	120 
    -- CP-element group 12: 	99 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	37 
    -- CP-element group 12: 	58 
    -- CP-element group 12: 	79 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	158 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	117 
    -- CP-element group 12: 	136 
    -- CP-element group 12: 	97 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	34 
    -- CP-element group 12: 	55 
    -- CP-element group 12: 	76 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1285_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1300_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1295_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1290_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1304_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1276_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1280_sample_completed_
      -- 
    outputPort_4_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(139) & outputPort_4_Daemon_CP_1900_elements(120) & outputPort_4_Daemon_CP_1900_elements(99) & outputPort_4_Daemon_CP_1900_elements(18) & outputPort_4_Daemon_CP_1900_elements(37) & outputPort_4_Daemon_CP_1900_elements(58) & outputPort_4_Daemon_CP_1900_elements(79);
      gj_outputPort_4_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	98 
    -- CP-element group 13: 	137 
    -- CP-element group 13: 	118 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	35 
    -- CP-element group 13: 	56 
    -- CP-element group 13: 	77 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	80 
    -- CP-element group 13: 	121 
    -- CP-element group 13: 	100 
    -- CP-element group 13: 	19 
    -- CP-element group 13: 	38 
    -- CP-element group 13: 	59 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1304_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/aggregated_phi_update_req
      -- 
    outputPort_4_Daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(98) & outputPort_4_Daemon_CP_1900_elements(137) & outputPort_4_Daemon_CP_1900_elements(118) & outputPort_4_Daemon_CP_1900_elements(16) & outputPort_4_Daemon_CP_1900_elements(35) & outputPort_4_Daemon_CP_1900_elements(56) & outputPort_4_Daemon_CP_1900_elements(77);
      gj_outputPort_4_Daemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	140 
    -- CP-element group 14: 	122 
    -- CP-element group 14: 	81 
    -- CP-element group 14: 	101 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	60 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/aggregated_phi_update_ack
      -- 
    outputPort_4_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(140) & outputPort_4_Daemon_CP_1900_elements(122) & outputPort_4_Daemon_CP_1900_elements(81) & outputPort_4_Daemon_CP_1900_elements(101) & outputPort_4_Daemon_CP_1900_elements(20) & outputPort_4_Daemon_CP_1900_elements(39) & outputPort_4_Daemon_CP_1900_elements(60);
      gj_outputPort_4_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1276_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	155 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1276_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(155);
      gj_outputPort_4_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1276_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(17) <= outputPort_4_Daemon_CP_1900_elements(11);
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1276_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1276_update_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(19) <= outputPort_4_Daemon_CP_1900_elements(13);
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	154 
    -- CP-element group 20: 	14 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1276_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1276_update_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1276_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(21) <= outputPort_4_Daemon_CP_1900_elements(7);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1276_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1276_loopback_sample_req_ps
      -- 
    phi_stmt_1276_loopback_sample_req_1939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1276_loopback_sample_req_1939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(22), ack => phi_stmt_1276_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1276_entry_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(23) <= outputPort_4_Daemon_CP_1900_elements(8);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1276_entry_sample_req
      -- CP-element group 24: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1276_entry_sample_req_ps
      -- 
    phi_stmt_1276_entry_sample_req_1942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1276_entry_sample_req_1942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(24), ack => phi_stmt_1276_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1276_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1276_phi_mux_ack_ps
      -- 
    phi_stmt_1276_phi_mux_ack_1945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1276_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_8_1278_sample_start__ps
      -- CP-element group 26: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_8_1278_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_8_1278_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_8_1278_sample_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_8_1278_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_8_1278_update_start_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_8_1278_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(28) <= outputPort_4_Daemon_CP_1900_elements(29);
    -- CP-element group 29:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	28 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_8_1278_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(29) is a control-delay.
    cp_element_29_delay: control_delay_element  generic map(name => " 29_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_1900_elements(27), ack => outputPort_4_Daemon_CP_1900_elements(29), clk => clk, reset =>reset);
    -- CP-element group 30:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_down_counter_1279_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_down_counter_1279_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_down_counter_1279_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_down_counter_1279_Sample/req
      -- 
    req_1966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(30), ack => next_down_counter_1387_1279_buf_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_down_counter_1279_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_down_counter_1279_update_start_
      -- CP-element group 31: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_down_counter_1279_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_down_counter_1279_Update/req
      -- 
    req_1971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(31), ack => next_down_counter_1387_1279_buf_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_down_counter_1279_sample_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_down_counter_1279_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_down_counter_1279_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_down_counter_1279_Sample/ack
      -- 
    ack_1967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_1387_1279_buf_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(32)); -- 
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_down_counter_1279_update_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_down_counter_1279_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_down_counter_1279_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_down_counter_1279_Update/ack
      -- 
    ack_1972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_1387_1279_buf_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(33)); -- 
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	9 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	12 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	11 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1280_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	155 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	13 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1280_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(155);
      gj_outputPort_4_Daemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	11 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1280_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(36) <= outputPort_4_Daemon_CP_1900_elements(11);
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	12 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1280_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1280_update_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(38) <= outputPort_4_Daemon_CP_1900_elements(13);
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	154 
    -- CP-element group 39: 	14 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1280_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1280_update_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	7 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1280_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(40) <= outputPort_4_Daemon_CP_1900_elements(7);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1280_loopback_sample_req
      -- CP-element group 41: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1280_loopback_sample_req_ps
      -- 
    phi_stmt_1280_loopback_sample_req_1983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1280_loopback_sample_req_1983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(41), ack => phi_stmt_1280_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	8 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1280_entry_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(42) <= outputPort_4_Daemon_CP_1900_elements(8);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1280_entry_sample_req
      -- CP-element group 43: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1280_entry_sample_req_ps
      -- 
    phi_stmt_1280_entry_sample_req_1986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1280_entry_sample_req_1986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(43), ack => phi_stmt_1280_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1280_phi_mux_ack_ps
      -- CP-element group 44: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1280_phi_mux_ack
      -- 
    phi_stmt_1280_phi_mux_ack_1989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1280_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1282_sample_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1282_sample_start__ps
      -- CP-element group 45: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1282_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1282_sample_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1282_update_start__ps
      -- CP-element group 46: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1282_update_start_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1282_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(47) <= outputPort_4_Daemon_CP_1900_elements(48);
    -- CP-element group 48:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	47 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1282_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(48) is a control-delay.
    cp_element_48_delay: control_delay_element  generic map(name => " 48_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_1900_elements(46), ack => outputPort_4_Daemon_CP_1900_elements(48), clk => clk, reset =>reset);
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_1_4_1284_sample_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_1_4_1284_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	54 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_1_4_1284_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_1_4_1284_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_1_4_1284_Sample/rr
      -- 
    rr_2010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(51), ack => RPIPE_noblock_obuf_1_4_1284_inst_req_0); -- 
    outputPort_4_Daemon_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(49) & outputPort_4_Daemon_CP_1900_elements(54);
      gj_outputPort_4_Daemon_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: 	53 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_1_4_1284_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_1_4_1284_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_1_4_1284_Update/cr
      -- 
    cr_2015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(52), ack => RPIPE_noblock_obuf_1_4_1284_inst_req_1); -- 
    outputPort_4_Daemon_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(50) & outputPort_4_Daemon_CP_1900_elements(53);
      gj_outputPort_4_Daemon_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	52 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_1_4_1284_sample_completed__ps
      -- CP-element group 53: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_1_4_1284_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_1_4_1284_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_1_4_1284_Sample/ra
      -- 
    ra_2011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_4_1284_inst_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(53)); -- 
    -- CP-element group 54:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	51 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_1_4_1284_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_1_4_1284_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_1_4_1284_update_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_1_4_1284_Update/$exit
      -- 
    ca_2016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_4_1284_inst_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(54)); -- 
    -- CP-element group 55:  join  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	9 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	12 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	11 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1285_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	9 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	155 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	13 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1285_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(155);
      gj_outputPort_4_Daemon_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	11 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1285_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(57) <= outputPort_4_Daemon_CP_1900_elements(11);
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	12 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1285_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	13 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1285_update_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(59) <= outputPort_4_Daemon_CP_1900_elements(13);
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	154 
    -- CP-element group 60: 	14 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1285_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1285_update_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	7 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1285_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(61) <= outputPort_4_Daemon_CP_1900_elements(7);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1285_loopback_sample_req_ps
      -- CP-element group 62: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1285_loopback_sample_req
      -- 
    phi_stmt_1285_loopback_sample_req_2027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1285_loopback_sample_req_2027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(62), ack => phi_stmt_1285_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	8 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1285_entry_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(63) <= outputPort_4_Daemon_CP_1900_elements(8);
    -- CP-element group 64:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1285_entry_sample_req_ps
      -- CP-element group 64: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1285_entry_sample_req
      -- 
    phi_stmt_1285_entry_sample_req_2030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1285_entry_sample_req_2030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(64), ack => phi_stmt_1285_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1285_phi_mux_ack_ps
      -- CP-element group 65: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1285_phi_mux_ack
      -- 
    phi_stmt_1285_phi_mux_ack_2033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1285_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(65)); -- 
    -- CP-element group 66:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1287_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1287_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1287_sample_completed__ps
      -- CP-element group 66: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1287_sample_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1287_update_start_
      -- CP-element group 67: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1287_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1287_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(68) <= outputPort_4_Daemon_CP_1900_elements(69);
    -- CP-element group 69:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	68 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1287_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(69) is a control-delay.
    cp_element_69_delay: control_delay_element  generic map(name => " 69_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_1900_elements(67), ack => outputPort_4_Daemon_CP_1900_elements(69), clk => clk, reset =>reset);
    -- CP-element group 70:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_2_4_1289_sample_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(70) is bound as output of CP function.
    -- CP-element group 71:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_2_4_1289_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: marked-predecessors 
    -- CP-element group 72: 	75 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_2_4_1289_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_2_4_1289_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_2_4_1289_Sample/rr
      -- 
    rr_2054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(72), ack => RPIPE_noblock_obuf_2_4_1289_inst_req_0); -- 
    outputPort_4_Daemon_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(70) & outputPort_4_Daemon_CP_1900_elements(75);
      gj_outputPort_4_Daemon_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: 	74 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_2_4_1289_update_start_
      -- CP-element group 73: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_2_4_1289_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_2_4_1289_Update/cr
      -- 
    cr_2059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(73), ack => RPIPE_noblock_obuf_2_4_1289_inst_req_1); -- 
    outputPort_4_Daemon_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(71) & outputPort_4_Daemon_CP_1900_elements(74);
      gj_outputPort_4_Daemon_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	73 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_2_4_1289_sample_completed__ps
      -- CP-element group 74: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_2_4_1289_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_2_4_1289_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_2_4_1289_Sample/ra
      -- 
    ra_2055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_4_1289_inst_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(74)); -- 
    -- CP-element group 75:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	72 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_2_4_1289_update_completed__ps
      -- CP-element group 75: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_2_4_1289_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_2_4_1289_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_2_4_1289_Update/ca
      -- 
    ca_2060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_4_1289_inst_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(75)); -- 
    -- CP-element group 76:  join  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	9 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	12 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	11 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1290_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	9 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	155 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	13 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1290_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(155);
      gj_outputPort_4_Daemon_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	11 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1290_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(78) <= outputPort_4_Daemon_CP_1900_elements(11);
    -- CP-element group 79:  join  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	12 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1290_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	13 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1290_update_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(80) <= outputPort_4_Daemon_CP_1900_elements(13);
    -- CP-element group 81:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	154 
    -- CP-element group 81: 	14 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1290_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1290_update_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	7 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1290_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(82) <= outputPort_4_Daemon_CP_1900_elements(7);
    -- CP-element group 83:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1290_loopback_sample_req_ps
      -- CP-element group 83: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1290_loopback_sample_req
      -- 
    phi_stmt_1290_loopback_sample_req_2071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1290_loopback_sample_req_2071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(83), ack => phi_stmt_1290_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(83) is bound as output of CP function.
    -- CP-element group 84:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	8 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1290_entry_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(84) <= outputPort_4_Daemon_CP_1900_elements(8);
    -- CP-element group 85:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1290_entry_sample_req
      -- CP-element group 85: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1290_entry_sample_req_ps
      -- 
    phi_stmt_1290_entry_sample_req_2074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1290_entry_sample_req_2074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(85), ack => phi_stmt_1290_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1290_phi_mux_ack_ps
      -- CP-element group 86: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1290_phi_mux_ack
      -- 
    phi_stmt_1290_phi_mux_ack_2077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1290_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(86)); -- 
    -- CP-element group 87:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1292_sample_completed__ps
      -- CP-element group 87: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1292_sample_start__ps
      -- CP-element group 87: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1292_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1292_sample_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1292_update_start__ps
      -- CP-element group 88: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1292_update_start_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	90 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1292_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(89) <= outputPort_4_Daemon_CP_1900_elements(90);
    -- CP-element group 90:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	89 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1292_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(90) is a control-delay.
    cp_element_90_delay: control_delay_element  generic map(name => " 90_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_1900_elements(88), ack => outputPort_4_Daemon_CP_1900_elements(90), clk => clk, reset =>reset);
    -- CP-element group 91:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_3_4_1294_sample_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(91) is bound as output of CP function.
    -- CP-element group 92:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_3_4_1294_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(92) is bound as output of CP function.
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	96 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_3_4_1294_Sample/rr
      -- CP-element group 93: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_3_4_1294_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_3_4_1294_sample_start_
      -- 
    rr_2098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(93), ack => RPIPE_noblock_obuf_3_4_1294_inst_req_0); -- 
    outputPort_4_Daemon_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(91) & outputPort_4_Daemon_CP_1900_elements(96);
      gj_outputPort_4_Daemon_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	95 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_3_4_1294_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_3_4_1294_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_3_4_1294_update_start_
      -- 
    cr_2103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(94), ack => RPIPE_noblock_obuf_3_4_1294_inst_req_1); -- 
    outputPort_4_Daemon_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(92) & outputPort_4_Daemon_CP_1900_elements(95);
      gj_outputPort_4_Daemon_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	94 
    -- CP-element group 95:  members (4) 
      -- CP-element group 95: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_3_4_1294_Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_3_4_1294_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_3_4_1294_sample_completed__ps
      -- CP-element group 95: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_3_4_1294_sample_completed_
      -- 
    ra_2099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_4_1294_inst_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(95)); -- 
    -- CP-element group 96:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	93 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_3_4_1294_Update/ca
      -- CP-element group 96: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_3_4_1294_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_3_4_1294_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_3_4_1294_update_completed__ps
      -- 
    ca_2104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_4_1294_inst_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(96)); -- 
    -- CP-element group 97:  join  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	9 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	12 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	11 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1295_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	9 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	155 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	13 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1295_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(155);
      gj_outputPort_4_Daemon_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  join  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	12 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1295_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(99) is bound as output of CP function.
    -- CP-element group 100:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	13 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1295_update_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(100) <= outputPort_4_Daemon_CP_1900_elements(13);
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	154 
    -- CP-element group 101: 	14 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1295_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1295_update_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(101) is bound as output of CP function.
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	7 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1295_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(102) <= outputPort_4_Daemon_CP_1900_elements(7);
    -- CP-element group 103:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1295_loopback_sample_req
      -- CP-element group 103: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1295_loopback_sample_req_ps
      -- 
    phi_stmt_1295_loopback_sample_req_2115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1295_loopback_sample_req_2115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(103), ack => phi_stmt_1295_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(103) is bound as output of CP function.
    -- CP-element group 104:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	8 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1295_entry_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(104) <= outputPort_4_Daemon_CP_1900_elements(8);
    -- CP-element group 105:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1295_entry_sample_req
      -- CP-element group 105: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1295_entry_sample_req_ps
      -- 
    phi_stmt_1295_entry_sample_req_2118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1295_entry_sample_req_2118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(105), ack => phi_stmt_1295_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(105) is bound as output of CP function.
    -- CP-element group 106:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1295_phi_mux_ack
      -- CP-element group 106: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1295_phi_mux_ack_ps
      -- 
    phi_stmt_1295_phi_mux_ack_2121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1295_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(106)); -- 
    -- CP-element group 107:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (4) 
      -- CP-element group 107: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1297_sample_start__ps
      -- CP-element group 107: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1297_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1297_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1297_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(107) is bound as output of CP function.
    -- CP-element group 108:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1297_update_start_
      -- CP-element group 108: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1297_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(108) is bound as output of CP function.
    -- CP-element group 109:  join  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	110 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1297_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(109) <= outputPort_4_Daemon_CP_1900_elements(110);
    -- CP-element group 110:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	109 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_33_1297_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(110) is a control-delay.
    cp_element_110_delay: control_delay_element  generic map(name => " 110_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_1900_elements(108), ack => outputPort_4_Daemon_CP_1900_elements(110), clk => clk, reset =>reset);
    -- CP-element group 111:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_4_4_1299_sample_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(111) is bound as output of CP function.
    -- CP-element group 112:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_4_4_1299_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(112) is bound as output of CP function.
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	116 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_4_4_1299_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_4_4_1299_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_4_4_1299_Sample/rr
      -- 
    rr_2142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(113), ack => RPIPE_noblock_obuf_4_4_1299_inst_req_0); -- 
    outputPort_4_Daemon_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(111) & outputPort_4_Daemon_CP_1900_elements(116);
      gj_outputPort_4_Daemon_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	115 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_4_4_1299_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_4_4_1299_update_start_
      -- CP-element group 114: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_4_4_1299_Update/cr
      -- 
    cr_2147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(114), ack => RPIPE_noblock_obuf_4_4_1299_inst_req_1); -- 
    outputPort_4_Daemon_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(115) & outputPort_4_Daemon_CP_1900_elements(112);
      gj_outputPort_4_Daemon_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	114 
    -- CP-element group 115:  members (4) 
      -- CP-element group 115: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_4_4_1299_sample_completed__ps
      -- CP-element group 115: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_4_4_1299_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_4_4_1299_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_4_4_1299_Sample/ra
      -- 
    ra_2143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_4_1299_inst_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(115)); -- 
    -- CP-element group 116:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: marked-successors 
    -- CP-element group 116: 	113 
    -- CP-element group 116:  members (4) 
      -- CP-element group 116: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_4_4_1299_update_completed__ps
      -- CP-element group 116: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_4_4_1299_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_4_4_1299_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/RPIPE_noblock_obuf_4_4_1299_Update/ca
      -- 
    ca_2148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_4_1299_inst_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(116)); -- 
    -- CP-element group 117:  join  transition  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	9 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	12 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	11 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1300_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	9 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	155 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	13 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1300_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(155);
      gj_outputPort_4_Daemon_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	11 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1300_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(119) <= outputPort_4_Daemon_CP_1900_elements(11);
    -- CP-element group 120:  join  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	12 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1300_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(120) is bound as output of CP function.
    -- CP-element group 121:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	13 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1300_update_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(121) <= outputPort_4_Daemon_CP_1900_elements(13);
    -- CP-element group 122:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	154 
    -- CP-element group 122: 	14 
    -- CP-element group 122:  members (2) 
      -- CP-element group 122: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1300_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1300_update_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(122) is bound as output of CP function.
    -- CP-element group 123:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	7 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1300_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(123) <= outputPort_4_Daemon_CP_1900_elements(7);
    -- CP-element group 124:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (2) 
      -- CP-element group 124: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1300_loopback_sample_req
      -- CP-element group 124: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1300_loopback_sample_req_ps
      -- 
    phi_stmt_1300_loopback_sample_req_2159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1300_loopback_sample_req_2159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(124), ack => phi_stmt_1300_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(124) is bound as output of CP function.
    -- CP-element group 125:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	8 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1300_entry_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(125) <= outputPort_4_Daemon_CP_1900_elements(8);
    -- CP-element group 126:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1300_entry_sample_req_ps
      -- CP-element group 126: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1300_entry_sample_req
      -- 
    phi_stmt_1300_entry_sample_req_2162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1300_entry_sample_req_2162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(126), ack => phi_stmt_1300_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(126) is bound as output of CP function.
    -- CP-element group 127:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1300_phi_mux_ack_ps
      -- CP-element group 127: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1300_phi_mux_ack
      -- 
    phi_stmt_1300_phi_mux_ack_2165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1300_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(127)); -- 
    -- CP-element group 128:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (4) 
      -- CP-element group 128: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_3_1302_sample_completed_
      -- CP-element group 128: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_3_1302_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_3_1302_sample_start__ps
      -- CP-element group 128: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_3_1302_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(128) is bound as output of CP function.
    -- CP-element group 129:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (2) 
      -- CP-element group 129: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_3_1302_update_start_
      -- CP-element group 129: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_3_1302_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(129) is bound as output of CP function.
    -- CP-element group 130:  join  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_3_1302_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(130) <= outputPort_4_Daemon_CP_1900_elements(131);
    -- CP-element group 131:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	130 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ZERO_3_1302_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(131) is a control-delay.
    cp_element_131_delay: control_delay_element  generic map(name => " 131_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_1900_elements(129), ack => outputPort_4_Daemon_CP_1900_elements(131), clk => clk, reset =>reset);
    -- CP-element group 132:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (4) 
      -- CP-element group 132: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_active_packet_1303_sample_start__ps
      -- CP-element group 132: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_active_packet_1303_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_active_packet_1303_Sample/req
      -- CP-element group 132: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_active_packet_1303_sample_start_
      -- 
    req_2186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(132), ack => next_active_packet_1367_1303_buf_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(132) is bound as output of CP function.
    -- CP-element group 133:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	135 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_active_packet_1303_update_start_
      -- CP-element group 133: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_active_packet_1303_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_active_packet_1303_update_start__ps
      -- CP-element group 133: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_active_packet_1303_Update/req
      -- 
    req_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(133), ack => next_active_packet_1367_1303_buf_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(133) is bound as output of CP function.
    -- CP-element group 134:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_active_packet_1303_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_active_packet_1303_Sample/$exit
      -- CP-element group 134: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_active_packet_1303_sample_completed__ps
      -- CP-element group 134: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_active_packet_1303_Sample/ack
      -- 
    ack_2187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_1367_1303_buf_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(134)); -- 
    -- CP-element group 135:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	133 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (4) 
      -- CP-element group 135: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_active_packet_1303_update_completed_
      -- CP-element group 135: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_active_packet_1303_Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_active_packet_1303_update_completed__ps
      -- CP-element group 135: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_active_packet_1303_Update/ack
      -- 
    ack_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_1367_1303_buf_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(135)); -- 
    -- CP-element group 136:  join  transition  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	9 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	12 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	11 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1304_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  join  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	9 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	155 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	13 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1304_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(155);
      gj_outputPort_4_Daemon_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	11 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1304_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(138) <= outputPort_4_Daemon_CP_1900_elements(11);
    -- CP-element group 139:  join  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	12 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1304_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(139) is bound as output of CP function.
    -- CP-element group 140:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	154 
    -- CP-element group 140: 	14 
    -- CP-element group 140:  members (2) 
      -- CP-element group 140: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1304_update_completed__ps
      -- CP-element group 140: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1304_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(140) is bound as output of CP function.
    -- CP-element group 141:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	7 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1304_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(141) <= outputPort_4_Daemon_CP_1900_elements(7);
    -- CP-element group 142:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1304_loopback_sample_req_ps
      -- CP-element group 142: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1304_loopback_sample_req
      -- 
    phi_stmt_1304_loopback_sample_req_2203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1304_loopback_sample_req_2203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(142), ack => phi_stmt_1304_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(142) is bound as output of CP function.
    -- CP-element group 143:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	8 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1304_entry_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(143) <= outputPort_4_Daemon_CP_1900_elements(8);
    -- CP-element group 144:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1304_entry_sample_req_ps
      -- CP-element group 144: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1304_entry_sample_req
      -- 
    phi_stmt_1304_entry_sample_req_2206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1304_entry_sample_req_2206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(144), ack => phi_stmt_1304_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1304_phi_mux_ack_ps
      -- CP-element group 145: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/phi_stmt_1304_phi_mux_ack
      -- 
    phi_stmt_1304_phi_mux_ack_2209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1304_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(145)); -- 
    -- CP-element group 146:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (4) 
      -- CP-element group 146: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ONE_3_1306_sample_completed_
      -- CP-element group 146: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ONE_3_1306_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ONE_3_1306_sample_completed__ps
      -- CP-element group 146: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ONE_3_1306_sample_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(146) is bound as output of CP function.
    -- CP-element group 147:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (2) 
      -- CP-element group 147: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ONE_3_1306_update_start__ps
      -- CP-element group 147: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ONE_3_1306_update_start_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(147) is bound as output of CP function.
    -- CP-element group 148:  join  transition  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	149 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (1) 
      -- CP-element group 148: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ONE_3_1306_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(148) <= outputPort_4_Daemon_CP_1900_elements(149);
    -- CP-element group 149:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	148 
    -- CP-element group 149:  members (1) 
      -- CP-element group 149: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_ONE_3_1306_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(149) is a control-delay.
    cp_element_149_delay: control_delay_element  generic map(name => " 149_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_1900_elements(147), ack => outputPort_4_Daemon_CP_1900_elements(149), clk => clk, reset =>reset);
    -- CP-element group 150:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (4) 
      -- CP-element group 150: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_pkt_priority_1307_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_pkt_priority_1307_Sample/req
      -- CP-element group 150: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_pkt_priority_1307_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_pkt_priority_1307_sample_start__ps
      -- 
    req_2230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(150), ack => next_pkt_priority_1367_1307_buf_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(150) is bound as output of CP function.
    -- CP-element group 151:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (4) 
      -- CP-element group 151: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_pkt_priority_1307_update_start__ps
      -- CP-element group 151: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_pkt_priority_1307_Update/req
      -- CP-element group 151: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_pkt_priority_1307_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_pkt_priority_1307_update_start_
      -- 
    req_2235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(151), ack => next_pkt_priority_1367_1307_buf_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(151) is bound as output of CP function.
    -- CP-element group 152:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (4) 
      -- CP-element group 152: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_pkt_priority_1307_Sample/ack
      -- CP-element group 152: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_pkt_priority_1307_sample_completed__ps
      -- CP-element group 152: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_pkt_priority_1307_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_pkt_priority_1307_sample_completed_
      -- 
    ack_2231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pkt_priority_1367_1307_buf_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(152)); -- 
    -- CP-element group 153:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (4) 
      -- CP-element group 153: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_pkt_priority_1307_Update/ack
      -- CP-element group 153: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_pkt_priority_1307_update_completed__ps
      -- CP-element group 153: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_pkt_priority_1307_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/R_next_pkt_priority_1307_update_completed_
      -- 
    ack_2236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pkt_priority_1367_1307_buf_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	140 
    -- CP-element group 154: 	122 
    -- CP-element group 154: 	81 
    -- CP-element group 154: 	101 
    -- CP-element group 154: 	20 
    -- CP-element group 154: 	39 
    -- CP-element group 154: 	60 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/WPIPE_out_data_4_1494_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/WPIPE_out_data_4_1494_Sample/req
      -- CP-element group 154: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/WPIPE_out_data_4_1494_Sample/$entry
      -- 
    req_2245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(154), ack => WPIPE_out_data_4_1494_inst_req_0); -- 
    outputPort_4_Daemon_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(140) & outputPort_4_Daemon_CP_1900_elements(122) & outputPort_4_Daemon_CP_1900_elements(81) & outputPort_4_Daemon_CP_1900_elements(101) & outputPort_4_Daemon_CP_1900_elements(20) & outputPort_4_Daemon_CP_1900_elements(39) & outputPort_4_Daemon_CP_1900_elements(60) & outputPort_4_Daemon_CP_1900_elements(156);
      gj_outputPort_4_Daemon_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	98 
    -- CP-element group 155: 	137 
    -- CP-element group 155: 	118 
    -- CP-element group 155: 	16 
    -- CP-element group 155: 	35 
    -- CP-element group 155: 	56 
    -- CP-element group 155: 	77 
    -- CP-element group 155:  members (6) 
      -- CP-element group 155: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/WPIPE_out_data_4_1494_Update/req
      -- CP-element group 155: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/WPIPE_out_data_4_1494_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/WPIPE_out_data_4_1494_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/WPIPE_out_data_4_1494_Sample/ack
      -- CP-element group 155: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/WPIPE_out_data_4_1494_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/WPIPE_out_data_4_1494_update_start_
      -- 
    ack_2246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_4_1494_inst_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(155)); -- 
    req_2250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(155), ack => WPIPE_out_data_4_1494_inst_req_1); -- 
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	154 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/WPIPE_out_data_4_1494_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/WPIPE_out_data_4_1494_Update/ack
      -- CP-element group 156: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/WPIPE_out_data_4_1494_update_completed_
      -- 
    ack_2251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_4_1494_inst_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(156)); -- 
    -- CP-element group 157:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	9 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	10 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(157) is a control-delay.
    cp_element_157_delay: control_delay_element  generic map(name => " 157_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_1900_elements(9), ack => outputPort_4_Daemon_CP_1900_elements(157), clk => clk, reset =>reset);
    -- CP-element group 158:  join  transition  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: 	12 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	6 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_1273/do_while_stmt_1274/do_while_stmt_1274_loop_body/$exit
      -- 
    outputPort_4_Daemon_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(156) & outputPort_4_Daemon_CP_1900_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	5 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (2) 
      -- CP-element group 159: 	 branch_block_stmt_1273/do_while_stmt_1274/loop_exit/$exit
      -- CP-element group 159: 	 branch_block_stmt_1273/do_while_stmt_1274/loop_exit/ack
      -- 
    ack_2256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1274_branch_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	5 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (2) 
      -- CP-element group 160: 	 branch_block_stmt_1273/do_while_stmt_1274/loop_taken/$exit
      -- CP-element group 160: 	 branch_block_stmt_1273/do_while_stmt_1274/loop_taken/ack
      -- 
    ack_2260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1274_branch_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(160)); -- 
    -- CP-element group 161:  transition  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	3 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	1 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_1273/do_while_stmt_1274/$exit
      -- 
    outputPort_4_Daemon_CP_1900_elements(161) <= outputPort_4_Daemon_CP_1900_elements(3);
    outputPort_4_Daemon_do_while_stmt_1274_terminator_2261: loop_terminator -- 
      generic map (name => " outputPort_4_Daemon_do_while_stmt_1274_terminator_2261", max_iterations_in_flight =>7) 
      port map(loop_body_exit => outputPort_4_Daemon_CP_1900_elements(6),loop_continue => outputPort_4_Daemon_CP_1900_elements(160),loop_terminate => outputPort_4_Daemon_CP_1900_elements(159),loop_back => outputPort_4_Daemon_CP_1900_elements(4),loop_exit => outputPort_4_Daemon_CP_1900_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1276_phi_seq_1973_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_1900_elements(23);
      outputPort_4_Daemon_CP_1900_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(26);
      outputPort_4_Daemon_CP_1900_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(28);
      outputPort_4_Daemon_CP_1900_elements(24) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_1900_elements(21);
      outputPort_4_Daemon_CP_1900_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(32);
      outputPort_4_Daemon_CP_1900_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(33);
      outputPort_4_Daemon_CP_1900_elements(22) <= phi_mux_reqs(1);
      phi_stmt_1276_phi_seq_1973 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1276_phi_seq_1973") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_1900_elements(17), 
          phi_sample_ack => outputPort_4_Daemon_CP_1900_elements(18), 
          phi_update_req => outputPort_4_Daemon_CP_1900_elements(19), 
          phi_update_ack => outputPort_4_Daemon_CP_1900_elements(20), 
          phi_mux_ack => outputPort_4_Daemon_CP_1900_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1280_phi_seq_2017_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_1900_elements(42);
      outputPort_4_Daemon_CP_1900_elements(45)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(45);
      outputPort_4_Daemon_CP_1900_elements(46)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(47);
      outputPort_4_Daemon_CP_1900_elements(43) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_1900_elements(40);
      outputPort_4_Daemon_CP_1900_elements(49)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(53);
      outputPort_4_Daemon_CP_1900_elements(50)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(54);
      outputPort_4_Daemon_CP_1900_elements(41) <= phi_mux_reqs(1);
      phi_stmt_1280_phi_seq_2017 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1280_phi_seq_2017") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_1900_elements(36), 
          phi_sample_ack => outputPort_4_Daemon_CP_1900_elements(37), 
          phi_update_req => outputPort_4_Daemon_CP_1900_elements(38), 
          phi_update_ack => outputPort_4_Daemon_CP_1900_elements(39), 
          phi_mux_ack => outputPort_4_Daemon_CP_1900_elements(44), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1285_phi_seq_2061_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_1900_elements(63);
      outputPort_4_Daemon_CP_1900_elements(66)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(66);
      outputPort_4_Daemon_CP_1900_elements(67)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(68);
      outputPort_4_Daemon_CP_1900_elements(64) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_1900_elements(61);
      outputPort_4_Daemon_CP_1900_elements(70)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(74);
      outputPort_4_Daemon_CP_1900_elements(71)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(75);
      outputPort_4_Daemon_CP_1900_elements(62) <= phi_mux_reqs(1);
      phi_stmt_1285_phi_seq_2061 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1285_phi_seq_2061") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_1900_elements(57), 
          phi_sample_ack => outputPort_4_Daemon_CP_1900_elements(58), 
          phi_update_req => outputPort_4_Daemon_CP_1900_elements(59), 
          phi_update_ack => outputPort_4_Daemon_CP_1900_elements(60), 
          phi_mux_ack => outputPort_4_Daemon_CP_1900_elements(65), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1290_phi_seq_2105_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_1900_elements(84);
      outputPort_4_Daemon_CP_1900_elements(87)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(87);
      outputPort_4_Daemon_CP_1900_elements(88)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(89);
      outputPort_4_Daemon_CP_1900_elements(85) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_1900_elements(82);
      outputPort_4_Daemon_CP_1900_elements(91)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(95);
      outputPort_4_Daemon_CP_1900_elements(92)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(96);
      outputPort_4_Daemon_CP_1900_elements(83) <= phi_mux_reqs(1);
      phi_stmt_1290_phi_seq_2105 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1290_phi_seq_2105") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_1900_elements(78), 
          phi_sample_ack => outputPort_4_Daemon_CP_1900_elements(79), 
          phi_update_req => outputPort_4_Daemon_CP_1900_elements(80), 
          phi_update_ack => outputPort_4_Daemon_CP_1900_elements(81), 
          phi_mux_ack => outputPort_4_Daemon_CP_1900_elements(86), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1295_phi_seq_2149_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_1900_elements(104);
      outputPort_4_Daemon_CP_1900_elements(107)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(107);
      outputPort_4_Daemon_CP_1900_elements(108)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(109);
      outputPort_4_Daemon_CP_1900_elements(105) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_1900_elements(102);
      outputPort_4_Daemon_CP_1900_elements(111)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(115);
      outputPort_4_Daemon_CP_1900_elements(112)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(116);
      outputPort_4_Daemon_CP_1900_elements(103) <= phi_mux_reqs(1);
      phi_stmt_1295_phi_seq_2149 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1295_phi_seq_2149") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_1900_elements(11), 
          phi_sample_ack => outputPort_4_Daemon_CP_1900_elements(99), 
          phi_update_req => outputPort_4_Daemon_CP_1900_elements(100), 
          phi_update_ack => outputPort_4_Daemon_CP_1900_elements(101), 
          phi_mux_ack => outputPort_4_Daemon_CP_1900_elements(106), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1300_phi_seq_2193_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_1900_elements(125);
      outputPort_4_Daemon_CP_1900_elements(128)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(128);
      outputPort_4_Daemon_CP_1900_elements(129)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(130);
      outputPort_4_Daemon_CP_1900_elements(126) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_1900_elements(123);
      outputPort_4_Daemon_CP_1900_elements(132)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(134);
      outputPort_4_Daemon_CP_1900_elements(133)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(135);
      outputPort_4_Daemon_CP_1900_elements(124) <= phi_mux_reqs(1);
      phi_stmt_1300_phi_seq_2193 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1300_phi_seq_2193") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_1900_elements(119), 
          phi_sample_ack => outputPort_4_Daemon_CP_1900_elements(120), 
          phi_update_req => outputPort_4_Daemon_CP_1900_elements(121), 
          phi_update_ack => outputPort_4_Daemon_CP_1900_elements(122), 
          phi_mux_ack => outputPort_4_Daemon_CP_1900_elements(127), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1304_phi_seq_2237_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_1900_elements(143);
      outputPort_4_Daemon_CP_1900_elements(146)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(146);
      outputPort_4_Daemon_CP_1900_elements(147)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(148);
      outputPort_4_Daemon_CP_1900_elements(144) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_1900_elements(141);
      outputPort_4_Daemon_CP_1900_elements(150)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(152);
      outputPort_4_Daemon_CP_1900_elements(151)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(153);
      outputPort_4_Daemon_CP_1900_elements(142) <= phi_mux_reqs(1);
      phi_stmt_1304_phi_seq_2237 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1304_phi_seq_2237") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_1900_elements(138), 
          phi_sample_ack => outputPort_4_Daemon_CP_1900_elements(139), 
          phi_update_req => outputPort_4_Daemon_CP_1900_elements(13), 
          phi_update_ack => outputPort_4_Daemon_CP_1900_elements(140), 
          phi_mux_ack => outputPort_4_Daemon_CP_1900_elements(145), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1925_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= outputPort_4_Daemon_CP_1900_elements(7);
        preds(1)  <= outputPort_4_Daemon_CP_1900_elements(8);
        entry_tmerge_1925 : transition_merge -- 
          generic map(name => " entry_tmerge_1925")
          port map (preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u3_u1_1332_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1338_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1345_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1351_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1393_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1401_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1409_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1417_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1434_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1441_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1449_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1456_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1467_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1473_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1480_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1486_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_1374_wire : std_logic_vector(0 downto 0);
    signal MUX_1335_wire : std_logic_vector(0 downto 0);
    signal MUX_1341_wire : std_logic_vector(0 downto 0);
    signal MUX_1348_wire : std_logic_vector(0 downto 0);
    signal MUX_1354_wire : std_logic_vector(0 downto 0);
    signal MUX_1385_wire : std_logic_vector(7 downto 0);
    signal MUX_1438_wire : std_logic_vector(31 downto 0);
    signal MUX_1445_wire : std_logic_vector(31 downto 0);
    signal MUX_1453_wire : std_logic_vector(31 downto 0);
    signal MUX_1460_wire : std_logic_vector(31 downto 0);
    signal MUX_1470_wire : std_logic_vector(0 downto 0);
    signal MUX_1476_wire : std_logic_vector(0 downto 0);
    signal MUX_1483_wire : std_logic_vector(0 downto 0);
    signal MUX_1489_wire : std_logic_vector(0 downto 0);
    signal NEQ_u3_u1_1371_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1390_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1398_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1406_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1414_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1342_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1355_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1477_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1490_wire : std_logic_vector(0 downto 0);
    signal OR_u32_u32_1446_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_1461_wire : std_logic_vector(31 downto 0);
    signal RPIPE_noblock_obuf_1_4_1284_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_2_4_1289_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_3_4_1294_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_4_4_1299_wire : std_logic_vector(32 downto 0);
    signal R_ONE_3_1306_wire_constant : std_logic_vector(2 downto 0);
    signal R_ZERO_33_1282_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1287_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1292_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1297_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_3_1302_wire_constant : std_logic_vector(2 downto 0);
    signal R_ZERO_8_1278_wire_constant : std_logic_vector(7 downto 0);
    signal SUB_u8_u8_1383_wire : std_logic_vector(7 downto 0);
    signal active_packet_1300 : std_logic_vector(2 downto 0);
    signal data_to_out_1463 : std_logic_vector(31 downto 0);
    signal down_counter_1276 : std_logic_vector(7 downto 0);
    signal konst_1311_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1316_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1321_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1326_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1331_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1334_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1337_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1340_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1344_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1347_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1350_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1353_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1370_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1373_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1379_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1382_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1392_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1400_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1408_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1416_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1433_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1437_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1440_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1444_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1448_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1452_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1455_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1459_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1466_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1469_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1472_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1475_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1479_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1482_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1485_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1488_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1498_wire_constant : std_logic_vector(0 downto 0);
    signal next_active_packet_1367 : std_logic_vector(2 downto 0);
    signal next_active_packet_1367_1303_buffered : std_logic_vector(2 downto 0);
    signal next_down_counter_1387 : std_logic_vector(7 downto 0);
    signal next_down_counter_1387_1279_buffered : std_logic_vector(7 downto 0);
    signal next_pkt_priority_1367 : std_logic_vector(2 downto 0);
    signal next_pkt_priority_1367_1307_buffered : std_logic_vector(2 downto 0);
    signal p1_valid_1313 : std_logic_vector(0 downto 0);
    signal p2_valid_1318 : std_logic_vector(0 downto 0);
    signal p3_valid_1323 : std_logic_vector(0 downto 0);
    signal p4_valid_1328 : std_logic_vector(0 downto 0);
    signal pkt_1_e_word_1280 : std_logic_vector(32 downto 0);
    signal pkt_2_e_word_1285 : std_logic_vector(32 downto 0);
    signal pkt_3_e_word_1290 : std_logic_vector(32 downto 0);
    signal pkt_4_e_word_1295 : std_logic_vector(32 downto 0);
    signal pkt_priority_1304 : std_logic_vector(2 downto 0);
    signal read_from_1_1395 : std_logic_vector(0 downto 0);
    signal read_from_2_1403 : std_logic_vector(0 downto 0);
    signal read_from_3_1411 : std_logic_vector(0 downto 0);
    signal read_from_4_1419 : std_logic_vector(0 downto 0);
    signal send_flag_1492 : std_logic_vector(0 downto 0);
    signal slice_1436_wire : std_logic_vector(31 downto 0);
    signal slice_1443_wire : std_logic_vector(31 downto 0);
    signal slice_1451_wire : std_logic_vector(31 downto 0);
    signal slice_1458_wire : std_logic_vector(31 downto 0);
    signal started_new_packet_1376 : std_logic_vector(0 downto 0);
    signal valid_active_pkt_word_read_1357 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_ONE_3_1306_wire_constant <= "001";
    R_ZERO_33_1282_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1287_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1292_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1297_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_3_1302_wire_constant <= "000";
    R_ZERO_8_1278_wire_constant <= "00000000";
    konst_1311_wire_constant <= "000000000000000000000000000100000";
    konst_1316_wire_constant <= "000000000000000000000000000100000";
    konst_1321_wire_constant <= "000000000000000000000000000100000";
    konst_1326_wire_constant <= "000000000000000000000000000100000";
    konst_1331_wire_constant <= "001";
    konst_1334_wire_constant <= "0";
    konst_1337_wire_constant <= "010";
    konst_1340_wire_constant <= "0";
    konst_1344_wire_constant <= "011";
    konst_1347_wire_constant <= "0";
    konst_1350_wire_constant <= "100";
    konst_1353_wire_constant <= "0";
    konst_1370_wire_constant <= "000";
    konst_1373_wire_constant <= "00000000";
    konst_1379_wire_constant <= "00111111";
    konst_1382_wire_constant <= "00000001";
    konst_1392_wire_constant <= "001";
    konst_1400_wire_constant <= "010";
    konst_1408_wire_constant <= "011";
    konst_1416_wire_constant <= "100";
    konst_1433_wire_constant <= "001";
    konst_1437_wire_constant <= "00000000000000000000000000000000";
    konst_1440_wire_constant <= "010";
    konst_1444_wire_constant <= "00000000000000000000000000000000";
    konst_1448_wire_constant <= "011";
    konst_1452_wire_constant <= "00000000000000000000000000000000";
    konst_1455_wire_constant <= "100";
    konst_1459_wire_constant <= "00000000000000000000000000000000";
    konst_1466_wire_constant <= "001";
    konst_1469_wire_constant <= "0";
    konst_1472_wire_constant <= "010";
    konst_1475_wire_constant <= "0";
    konst_1479_wire_constant <= "011";
    konst_1482_wire_constant <= "0";
    konst_1485_wire_constant <= "100";
    konst_1488_wire_constant <= "0";
    konst_1498_wire_constant <= "1";
    phi_stmt_1276: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_8_1278_wire_constant & next_down_counter_1387_1279_buffered;
      req <= phi_stmt_1276_req_0 & phi_stmt_1276_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1276",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1276_ack_0,
          idata => idata,
          odata => down_counter_1276,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1276
    phi_stmt_1280: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1282_wire_constant & RPIPE_noblock_obuf_1_4_1284_wire;
      req <= phi_stmt_1280_req_0 & phi_stmt_1280_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1280",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1280_ack_0,
          idata => idata,
          odata => pkt_1_e_word_1280,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1280
    phi_stmt_1285: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1287_wire_constant & RPIPE_noblock_obuf_2_4_1289_wire;
      req <= phi_stmt_1285_req_0 & phi_stmt_1285_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1285",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1285_ack_0,
          idata => idata,
          odata => pkt_2_e_word_1285,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1285
    phi_stmt_1290: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1292_wire_constant & RPIPE_noblock_obuf_3_4_1294_wire;
      req <= phi_stmt_1290_req_0 & phi_stmt_1290_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1290",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1290_ack_0,
          idata => idata,
          odata => pkt_3_e_word_1290,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1290
    phi_stmt_1295: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1297_wire_constant & RPIPE_noblock_obuf_4_4_1299_wire;
      req <= phi_stmt_1295_req_0 & phi_stmt_1295_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1295",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1295_ack_0,
          idata => idata,
          odata => pkt_4_e_word_1295,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1295
    phi_stmt_1300: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_3_1302_wire_constant & next_active_packet_1367_1303_buffered;
      req <= phi_stmt_1300_req_0 & phi_stmt_1300_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1300",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1300_ack_0,
          idata => idata,
          odata => active_packet_1300,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1300
    phi_stmt_1304: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ONE_3_1306_wire_constant & next_pkt_priority_1367_1307_buffered;
      req <= phi_stmt_1304_req_0 & phi_stmt_1304_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1304",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1304_ack_0,
          idata => idata,
          odata => pkt_priority_1304,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1304
    -- flow-through select operator MUX_1335_inst
    MUX_1335_wire <= p1_valid_1313 when (EQ_u3_u1_1332_wire(0) /=  '0') else konst_1334_wire_constant;
    -- flow-through select operator MUX_1341_inst
    MUX_1341_wire <= p2_valid_1318 when (EQ_u3_u1_1338_wire(0) /=  '0') else konst_1340_wire_constant;
    -- flow-through select operator MUX_1348_inst
    MUX_1348_wire <= p3_valid_1323 when (EQ_u3_u1_1345_wire(0) /=  '0') else konst_1347_wire_constant;
    -- flow-through select operator MUX_1354_inst
    MUX_1354_wire <= p4_valid_1328 when (EQ_u3_u1_1351_wire(0) /=  '0') else konst_1353_wire_constant;
    -- flow-through select operator MUX_1385_inst
    MUX_1385_wire <= SUB_u8_u8_1383_wire when (valid_active_pkt_word_read_1357(0) /=  '0') else down_counter_1276;
    -- flow-through select operator MUX_1386_inst
    next_down_counter_1387 <= konst_1379_wire_constant when (started_new_packet_1376(0) /=  '0') else MUX_1385_wire;
    -- flow-through select operator MUX_1438_inst
    MUX_1438_wire <= slice_1436_wire when (EQ_u3_u1_1434_wire(0) /=  '0') else konst_1437_wire_constant;
    -- flow-through select operator MUX_1445_inst
    MUX_1445_wire <= slice_1443_wire when (EQ_u3_u1_1441_wire(0) /=  '0') else konst_1444_wire_constant;
    -- flow-through select operator MUX_1453_inst
    MUX_1453_wire <= slice_1451_wire when (EQ_u3_u1_1449_wire(0) /=  '0') else konst_1452_wire_constant;
    -- flow-through select operator MUX_1460_inst
    MUX_1460_wire <= slice_1458_wire when (EQ_u3_u1_1456_wire(0) /=  '0') else konst_1459_wire_constant;
    -- flow-through select operator MUX_1470_inst
    MUX_1470_wire <= p1_valid_1313 when (EQ_u3_u1_1467_wire(0) /=  '0') else konst_1469_wire_constant;
    -- flow-through select operator MUX_1476_inst
    MUX_1476_wire <= p2_valid_1318 when (EQ_u3_u1_1473_wire(0) /=  '0') else konst_1475_wire_constant;
    -- flow-through select operator MUX_1483_inst
    MUX_1483_wire <= p3_valid_1323 when (EQ_u3_u1_1480_wire(0) /=  '0') else konst_1482_wire_constant;
    -- flow-through select operator MUX_1489_inst
    MUX_1489_wire <= p4_valid_1328 when (EQ_u3_u1_1486_wire(0) /=  '0') else konst_1488_wire_constant;
    -- flow-through slice operator slice_1436_inst
    slice_1436_wire <= pkt_1_e_word_1280(31 downto 0);
    -- flow-through slice operator slice_1443_inst
    slice_1443_wire <= pkt_2_e_word_1285(31 downto 0);
    -- flow-through slice operator slice_1451_inst
    slice_1451_wire <= pkt_3_e_word_1290(31 downto 0);
    -- flow-through slice operator slice_1458_inst
    slice_1458_wire <= pkt_4_e_word_1295(31 downto 0);
    next_active_packet_1367_1303_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_active_packet_1367_1303_buf_req_0;
      next_active_packet_1367_1303_buf_ack_0<= wack(0);
      rreq(0) <= next_active_packet_1367_1303_buf_req_1;
      next_active_packet_1367_1303_buf_ack_1<= rack(0);
      next_active_packet_1367_1303_buf : InterlockBuffer generic map ( -- 
        name => "next_active_packet_1367_1303_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_active_packet_1367,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_active_packet_1367_1303_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_down_counter_1387_1279_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_down_counter_1387_1279_buf_req_0;
      next_down_counter_1387_1279_buf_ack_0<= wack(0);
      rreq(0) <= next_down_counter_1387_1279_buf_req_1;
      next_down_counter_1387_1279_buf_ack_1<= rack(0);
      next_down_counter_1387_1279_buf : InterlockBuffer generic map ( -- 
        name => "next_down_counter_1387_1279_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_down_counter_1387,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_down_counter_1387_1279_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_pkt_priority_1367_1307_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_pkt_priority_1367_1307_buf_req_0;
      next_pkt_priority_1367_1307_buf_ack_0<= wack(0);
      rreq(0) <= next_pkt_priority_1367_1307_buf_req_1;
      next_pkt_priority_1367_1307_buf_ack_1<= rack(0);
      next_pkt_priority_1367_1307_buf : InterlockBuffer generic map ( -- 
        name => "next_pkt_priority_1367_1307_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_pkt_priority_1367,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_pkt_priority_1367_1307_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1274_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1498_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1274_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1274_branch_req_0,
          ack0 => do_while_stmt_1274_branch_ack_0,
          ack1 => do_while_stmt_1274_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator AND_u1_u1_1375_inst
    process(NEQ_u3_u1_1371_wire, EQ_u8_u1_1374_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NEQ_u3_u1_1371_wire, EQ_u8_u1_1374_wire, tmp_var);
      started_new_packet_1376 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_1312_inst
    process(pkt_1_e_word_1280) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_1_e_word_1280, konst_1311_wire_constant, tmp_var);
      p1_valid_1313 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_1317_inst
    process(pkt_2_e_word_1285) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_2_e_word_1285, konst_1316_wire_constant, tmp_var);
      p2_valid_1318 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_1322_inst
    process(pkt_3_e_word_1290) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_3_e_word_1290, konst_1321_wire_constant, tmp_var);
      p3_valid_1323 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_1327_inst
    process(pkt_4_e_word_1295) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_4_e_word_1295, konst_1326_wire_constant, tmp_var);
      p4_valid_1328 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1332_inst
    process(active_packet_1300) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1300, konst_1331_wire_constant, tmp_var);
      EQ_u3_u1_1332_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1338_inst
    process(active_packet_1300) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1300, konst_1337_wire_constant, tmp_var);
      EQ_u3_u1_1338_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1345_inst
    process(active_packet_1300) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1300, konst_1344_wire_constant, tmp_var);
      EQ_u3_u1_1345_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1351_inst
    process(active_packet_1300) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1300, konst_1350_wire_constant, tmp_var);
      EQ_u3_u1_1351_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1393_inst
    process(next_active_packet_1367) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1367, konst_1392_wire_constant, tmp_var);
      EQ_u3_u1_1393_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1401_inst
    process(next_active_packet_1367) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1367, konst_1400_wire_constant, tmp_var);
      EQ_u3_u1_1401_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1409_inst
    process(next_active_packet_1367) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1367, konst_1408_wire_constant, tmp_var);
      EQ_u3_u1_1409_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1417_inst
    process(next_active_packet_1367) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1367, konst_1416_wire_constant, tmp_var);
      EQ_u3_u1_1417_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1434_inst
    process(next_active_packet_1367) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1367, konst_1433_wire_constant, tmp_var);
      EQ_u3_u1_1434_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1441_inst
    process(next_active_packet_1367) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1367, konst_1440_wire_constant, tmp_var);
      EQ_u3_u1_1441_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1449_inst
    process(next_active_packet_1367) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1367, konst_1448_wire_constant, tmp_var);
      EQ_u3_u1_1449_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1456_inst
    process(next_active_packet_1367) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1367, konst_1455_wire_constant, tmp_var);
      EQ_u3_u1_1456_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1467_inst
    process(next_active_packet_1367) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1367, konst_1466_wire_constant, tmp_var);
      EQ_u3_u1_1467_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1473_inst
    process(next_active_packet_1367) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1367, konst_1472_wire_constant, tmp_var);
      EQ_u3_u1_1473_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1480_inst
    process(next_active_packet_1367) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1367, konst_1479_wire_constant, tmp_var);
      EQ_u3_u1_1480_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1486_inst
    process(next_active_packet_1367) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1367, konst_1485_wire_constant, tmp_var);
      EQ_u3_u1_1486_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_1374_inst
    process(down_counter_1276) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(down_counter_1276, konst_1373_wire_constant, tmp_var);
      EQ_u8_u1_1374_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u3_u1_1371_inst
    process(next_active_packet_1367) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(next_active_packet_1367, konst_1370_wire_constant, tmp_var);
      NEQ_u3_u1_1371_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1390_inst
    process(p1_valid_1313) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_1313, tmp_var);
      NOT_u1_u1_1390_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1398_inst
    process(p2_valid_1318) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_1318, tmp_var);
      NOT_u1_u1_1398_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1406_inst
    process(p3_valid_1323) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_1323, tmp_var);
      NOT_u1_u1_1406_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1414_inst
    process(p4_valid_1328) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_1328, tmp_var);
      NOT_u1_u1_1414_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1342_inst
    process(MUX_1335_wire, MUX_1341_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1335_wire, MUX_1341_wire, tmp_var);
      OR_u1_u1_1342_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1355_inst
    process(MUX_1348_wire, MUX_1354_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1348_wire, MUX_1354_wire, tmp_var);
      OR_u1_u1_1355_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1356_inst
    process(OR_u1_u1_1342_wire, OR_u1_u1_1355_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1342_wire, OR_u1_u1_1355_wire, tmp_var);
      valid_active_pkt_word_read_1357 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1394_inst
    process(NOT_u1_u1_1390_wire, EQ_u3_u1_1393_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1390_wire, EQ_u3_u1_1393_wire, tmp_var);
      read_from_1_1395 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1402_inst
    process(NOT_u1_u1_1398_wire, EQ_u3_u1_1401_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1398_wire, EQ_u3_u1_1401_wire, tmp_var);
      read_from_2_1403 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1410_inst
    process(NOT_u1_u1_1406_wire, EQ_u3_u1_1409_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1406_wire, EQ_u3_u1_1409_wire, tmp_var);
      read_from_3_1411 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1418_inst
    process(NOT_u1_u1_1414_wire, EQ_u3_u1_1417_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1414_wire, EQ_u3_u1_1417_wire, tmp_var);
      read_from_4_1419 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1477_inst
    process(MUX_1470_wire, MUX_1476_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1470_wire, MUX_1476_wire, tmp_var);
      OR_u1_u1_1477_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1490_inst
    process(MUX_1483_wire, MUX_1489_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1483_wire, MUX_1489_wire, tmp_var);
      OR_u1_u1_1490_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1491_inst
    process(OR_u1_u1_1477_wire, OR_u1_u1_1490_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1477_wire, OR_u1_u1_1490_wire, tmp_var);
      send_flag_1492 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1446_inst
    process(MUX_1438_wire, MUX_1445_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1438_wire, MUX_1445_wire, tmp_var);
      OR_u32_u32_1446_wire <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1461_inst
    process(MUX_1453_wire, MUX_1460_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1453_wire, MUX_1460_wire, tmp_var);
      OR_u32_u32_1461_wire <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1462_inst
    process(OR_u32_u32_1446_wire, OR_u32_u32_1461_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u32_u32_1446_wire, OR_u32_u32_1461_wire, tmp_var);
      data_to_out_1463 <= tmp_var; --
    end process;
    -- binary operator SUB_u8_u8_1383_inst
    process(down_counter_1276) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSub_proc(down_counter_1276, konst_1382_wire_constant, tmp_var);
      SUB_u8_u8_1383_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_noblock_obuf_1_4_1284_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_1_4_1284_inst_req_0;
      RPIPE_noblock_obuf_1_4_1284_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_1_4_1284_inst_req_1;
      RPIPE_noblock_obuf_1_4_1284_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_1_1395(0);
      RPIPE_noblock_obuf_1_4_1284_wire <= data_out(32 downto 0);
      noblock_obuf_1_4_read_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_4_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_4_read_0: InputPortRevised -- 
        generic map ( name => "noblock_obuf_1_4_read_0", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_1_4_pipe_read_req(0),
          oack => noblock_obuf_1_4_pipe_read_ack(0),
          odata => noblock_obuf_1_4_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_noblock_obuf_2_4_1289_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_2_4_1289_inst_req_0;
      RPIPE_noblock_obuf_2_4_1289_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_2_4_1289_inst_req_1;
      RPIPE_noblock_obuf_2_4_1289_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_2_1403(0);
      RPIPE_noblock_obuf_2_4_1289_wire <= data_out(32 downto 0);
      noblock_obuf_2_4_read_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_4_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_4_read_1: InputPortRevised -- 
        generic map ( name => "noblock_obuf_2_4_read_1", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_2_4_pipe_read_req(0),
          oack => noblock_obuf_2_4_pipe_read_ack(0),
          odata => noblock_obuf_2_4_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_noblock_obuf_3_4_1294_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_3_4_1294_inst_req_0;
      RPIPE_noblock_obuf_3_4_1294_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_3_4_1294_inst_req_1;
      RPIPE_noblock_obuf_3_4_1294_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_3_1411(0);
      RPIPE_noblock_obuf_3_4_1294_wire <= data_out(32 downto 0);
      noblock_obuf_3_4_read_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_4_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_4_read_2: InputPortRevised -- 
        generic map ( name => "noblock_obuf_3_4_read_2", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_3_4_pipe_read_req(0),
          oack => noblock_obuf_3_4_pipe_read_ack(0),
          odata => noblock_obuf_3_4_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_noblock_obuf_4_4_1299_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_4_4_1299_inst_req_0;
      RPIPE_noblock_obuf_4_4_1299_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_4_4_1299_inst_req_1;
      RPIPE_noblock_obuf_4_4_1299_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_4_1419(0);
      RPIPE_noblock_obuf_4_4_1299_wire <= data_out(32 downto 0);
      noblock_obuf_4_4_read_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_4_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_4_read_3: InputPortRevised -- 
        generic map ( name => "noblock_obuf_4_4_read_3", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_4_4_pipe_read_req(0),
          oack => noblock_obuf_4_4_pipe_read_ack(0),
          odata => noblock_obuf_4_4_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_out_data_4_1494_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_out_data_4_1494_inst_req_0;
      WPIPE_out_data_4_1494_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_out_data_4_1494_inst_req_1;
      WPIPE_out_data_4_1494_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_flag_1492(0);
      data_in <= data_to_out_1463;
      out_data_4_write_0_gI: SplitGuardInterface generic map(name => "out_data_4_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      out_data_4_write_0: OutputPortRevised -- 
        generic map ( name => "out_data_4", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => out_data_4_pipe_write_req(0),
          oack => out_data_4_pipe_write_ack(0),
          odata => out_data_4_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    volatile_operator_prioritySelect_3683: prioritySelect_Volatile port map(down_counter => down_counter_1276, active_packet => active_packet_1300, pkt_priority => pkt_priority_1304, p1_valid => p1_valid_1313, p2_valid => p2_valid_1318, p3_valid => p3_valid_1323, p4_valid => p4_valid_1328, next_active_packet => next_active_packet_1367, next_pkt_priority => next_pkt_priority_1367); 
    -- 
  end Block; -- data_path
  -- 
end outputPort_4_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity prioritySelect_Volatile is -- 
  port ( -- 
    down_counter : in  std_logic_vector(7 downto 0);
    active_packet : in  std_logic_vector(2 downto 0);
    pkt_priority : in  std_logic_vector(2 downto 0);
    p1_valid : in  std_logic_vector(0 downto 0);
    p2_valid : in  std_logic_vector(0 downto 0);
    p3_valid : in  std_logic_vector(0 downto 0);
    p4_valid : in  std_logic_vector(0 downto 0);
    next_active_packet : out  std_logic_vector(2 downto 0);
    next_pkt_priority : out  std_logic_vector(2 downto 0)-- 
  );
  -- 
end entity prioritySelect_Volatile;
architecture prioritySelect_Volatile_arch of prioritySelect_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(18-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal down_counter_buffer :  std_logic_vector(7 downto 0);
  signal active_packet_buffer :  std_logic_vector(2 downto 0);
  signal pkt_priority_buffer :  std_logic_vector(2 downto 0);
  signal p1_valid_buffer :  std_logic_vector(0 downto 0);
  signal p2_valid_buffer :  std_logic_vector(0 downto 0);
  signal p3_valid_buffer :  std_logic_vector(0 downto 0);
  signal p4_valid_buffer :  std_logic_vector(0 downto 0);
  -- output port buffer signals
  signal next_active_packet_buffer :  std_logic_vector(2 downto 0);
  signal next_pkt_priority_buffer :  std_logic_vector(2 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  down_counter_buffer <= down_counter;
  active_packet_buffer <= active_packet;
  pkt_priority_buffer <= pkt_priority;
  p1_valid_buffer <= p1_valid;
  p2_valid_buffer <= p2_valid;
  p3_valid_buffer <= p3_valid;
  p4_valid_buffer <= p4_valid;
  -- output handling  -------------------------------------------------------
  next_active_packet <= next_active_packet_buffer;
  next_pkt_priority <= next_pkt_priority_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_446_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_454_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_457_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_464_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_472_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_475_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_482_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_490_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_493_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_500_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_508_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_511_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_544_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_549_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_550_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_449_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_467_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_485_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_503_wire : std_logic_vector(0 downto 0);
    signal MUX_520_wire : std_logic_vector(2 downto 0);
    signal MUX_524_wire : std_logic_vector(2 downto 0);
    signal MUX_529_wire : std_logic_vector(2 downto 0);
    signal MUX_534_wire : std_logic_vector(2 downto 0);
    signal MUX_538_wire : std_logic_vector(2 downto 0);
    signal MUX_553_wire : std_logic_vector(2 downto 0);
    signal MUX_562_wire : std_logic_vector(2 downto 0);
    signal MUX_566_wire : std_logic_vector(2 downto 0);
    signal MUX_571_wire : std_logic_vector(2 downto 0);
    signal MUX_576_wire : std_logic_vector(2 downto 0);
    signal MUX_580_wire : std_logic_vector(2 downto 0);
    signal NOT_u1_u1_451_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_453_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_456_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_469_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_471_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_474_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_487_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_489_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_492_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_505_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_507_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_510_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_517_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_541_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_543_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_546_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_548_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_559_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_458_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_476_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_494_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_512_wire : std_logic_vector(0 downto 0);
    signal OR_u3_u3_525_wire : std_logic_vector(2 downto 0);
    signal OR_u3_u3_530_wire : std_logic_vector(2 downto 0);
    signal OR_u3_u3_539_wire : std_logic_vector(2 downto 0);
    signal OR_u3_u3_554_wire : std_logic_vector(2 downto 0);
    signal OR_u3_u3_567_wire : std_logic_vector(2 downto 0);
    signal OR_u3_u3_572_wire : std_logic_vector(2 downto 0);
    signal OR_u3_u3_581_wire : std_logic_vector(2 downto 0);
    signal d0_442 : std_logic_vector(0 downto 0);
    signal konst_440_wire_constant : std_logic_vector(7 downto 0);
    signal konst_448_wire_constant : std_logic_vector(2 downto 0);
    signal konst_466_wire_constant : std_logic_vector(2 downto 0);
    signal konst_484_wire_constant : std_logic_vector(2 downto 0);
    signal konst_502_wire_constant : std_logic_vector(2 downto 0);
    signal konst_519_wire_constant : std_logic_vector(2 downto 0);
    signal konst_522_wire_constant : std_logic_vector(2 downto 0);
    signal konst_523_wire_constant : std_logic_vector(2 downto 0);
    signal konst_527_wire_constant : std_logic_vector(2 downto 0);
    signal konst_528_wire_constant : std_logic_vector(2 downto 0);
    signal konst_532_wire_constant : std_logic_vector(2 downto 0);
    signal konst_533_wire_constant : std_logic_vector(2 downto 0);
    signal konst_536_wire_constant : std_logic_vector(2 downto 0);
    signal konst_537_wire_constant : std_logic_vector(2 downto 0);
    signal konst_552_wire_constant : std_logic_vector(2 downto 0);
    signal konst_561_wire_constant : std_logic_vector(2 downto 0);
    signal konst_564_wire_constant : std_logic_vector(2 downto 0);
    signal konst_565_wire_constant : std_logic_vector(2 downto 0);
    signal konst_569_wire_constant : std_logic_vector(2 downto 0);
    signal konst_570_wire_constant : std_logic_vector(2 downto 0);
    signal konst_574_wire_constant : std_logic_vector(2 downto 0);
    signal konst_575_wire_constant : std_logic_vector(2 downto 0);
    signal konst_578_wire_constant : std_logic_vector(2 downto 0);
    signal konst_579_wire_constant : std_logic_vector(2 downto 0);
    signal select_1_460 : std_logic_vector(0 downto 0);
    signal select_2_478 : std_logic_vector(0 downto 0);
    signal select_3_496 : std_logic_vector(0 downto 0);
    signal select_4_514 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    konst_440_wire_constant <= "00000000";
    konst_448_wire_constant <= "001";
    konst_466_wire_constant <= "010";
    konst_484_wire_constant <= "011";
    konst_502_wire_constant <= "100";
    konst_519_wire_constant <= "000";
    konst_522_wire_constant <= "001";
    konst_523_wire_constant <= "000";
    konst_527_wire_constant <= "010";
    konst_528_wire_constant <= "000";
    konst_532_wire_constant <= "011";
    konst_533_wire_constant <= "000";
    konst_536_wire_constant <= "100";
    konst_537_wire_constant <= "000";
    konst_552_wire_constant <= "000";
    konst_561_wire_constant <= "000";
    konst_564_wire_constant <= "010";
    konst_565_wire_constant <= "000";
    konst_569_wire_constant <= "011";
    konst_570_wire_constant <= "000";
    konst_574_wire_constant <= "100";
    konst_575_wire_constant <= "000";
    konst_578_wire_constant <= "001";
    konst_579_wire_constant <= "000";
    -- flow-through select operator MUX_520_inst
    MUX_520_wire <= active_packet_buffer when (NOT_u1_u1_517_wire(0) /=  '0') else konst_519_wire_constant;
    -- flow-through select operator MUX_524_inst
    MUX_524_wire <= konst_522_wire_constant when (select_1_460(0) /=  '0') else konst_523_wire_constant;
    -- flow-through select operator MUX_529_inst
    MUX_529_wire <= konst_527_wire_constant when (select_2_478(0) /=  '0') else konst_528_wire_constant;
    -- flow-through select operator MUX_534_inst
    MUX_534_wire <= konst_532_wire_constant when (select_3_496(0) /=  '0') else konst_533_wire_constant;
    -- flow-through select operator MUX_538_inst
    MUX_538_wire <= konst_536_wire_constant when (select_4_514(0) /=  '0') else konst_537_wire_constant;
    -- flow-through select operator MUX_553_inst
    MUX_553_wire <= active_packet_buffer when (AND_u1_u1_550_wire(0) /=  '0') else konst_552_wire_constant;
    -- flow-through select operator MUX_562_inst
    MUX_562_wire <= active_packet_buffer when (NOT_u1_u1_559_wire(0) /=  '0') else konst_561_wire_constant;
    -- flow-through select operator MUX_566_inst
    MUX_566_wire <= konst_564_wire_constant when (select_1_460(0) /=  '0') else konst_565_wire_constant;
    -- flow-through select operator MUX_571_inst
    MUX_571_wire <= konst_569_wire_constant when (select_2_478(0) /=  '0') else konst_570_wire_constant;
    -- flow-through select operator MUX_576_inst
    MUX_576_wire <= konst_574_wire_constant when (select_3_496(0) /=  '0') else konst_575_wire_constant;
    -- flow-through select operator MUX_580_inst
    MUX_580_wire <= konst_578_wire_constant when (select_4_514(0) /=  '0') else konst_579_wire_constant;
    -- binary operator AND_u1_u1_446_inst
    process(d0_442, p1_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(d0_442, p1_valid_buffer, tmp_var);
      AND_u1_u1_446_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_454_inst
    process(NOT_u1_u1_451_wire, NOT_u1_u1_453_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_451_wire, NOT_u1_u1_453_wire, tmp_var);
      AND_u1_u1_454_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_457_inst
    process(AND_u1_u1_454_wire, NOT_u1_u1_456_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_454_wire, NOT_u1_u1_456_wire, tmp_var);
      AND_u1_u1_457_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_459_inst
    process(AND_u1_u1_446_wire, OR_u1_u1_458_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_446_wire, OR_u1_u1_458_wire, tmp_var);
      select_1_460 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_464_inst
    process(d0_442, p2_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(d0_442, p2_valid_buffer, tmp_var);
      AND_u1_u1_464_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_472_inst
    process(NOT_u1_u1_469_wire, NOT_u1_u1_471_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_469_wire, NOT_u1_u1_471_wire, tmp_var);
      AND_u1_u1_472_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_475_inst
    process(AND_u1_u1_472_wire, NOT_u1_u1_474_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_472_wire, NOT_u1_u1_474_wire, tmp_var);
      AND_u1_u1_475_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_477_inst
    process(AND_u1_u1_464_wire, OR_u1_u1_476_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_464_wire, OR_u1_u1_476_wire, tmp_var);
      select_2_478 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_482_inst
    process(d0_442, p3_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(d0_442, p3_valid_buffer, tmp_var);
      AND_u1_u1_482_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_490_inst
    process(NOT_u1_u1_487_wire, NOT_u1_u1_489_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_487_wire, NOT_u1_u1_489_wire, tmp_var);
      AND_u1_u1_490_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_493_inst
    process(AND_u1_u1_490_wire, NOT_u1_u1_492_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_490_wire, NOT_u1_u1_492_wire, tmp_var);
      AND_u1_u1_493_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_495_inst
    process(AND_u1_u1_482_wire, OR_u1_u1_494_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_482_wire, OR_u1_u1_494_wire, tmp_var);
      select_3_496 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_500_inst
    process(d0_442, p4_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(d0_442, p4_valid_buffer, tmp_var);
      AND_u1_u1_500_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_508_inst
    process(NOT_u1_u1_505_wire, NOT_u1_u1_507_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_505_wire, NOT_u1_u1_507_wire, tmp_var);
      AND_u1_u1_508_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_511_inst
    process(AND_u1_u1_508_wire, NOT_u1_u1_510_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_508_wire, NOT_u1_u1_510_wire, tmp_var);
      AND_u1_u1_511_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_513_inst
    process(AND_u1_u1_500_wire, OR_u1_u1_512_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_500_wire, OR_u1_u1_512_wire, tmp_var);
      select_4_514 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_544_inst
    process(NOT_u1_u1_541_wire, NOT_u1_u1_543_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_541_wire, NOT_u1_u1_543_wire, tmp_var);
      AND_u1_u1_544_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_549_inst
    process(NOT_u1_u1_546_wire, NOT_u1_u1_548_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_546_wire, NOT_u1_u1_548_wire, tmp_var);
      AND_u1_u1_549_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_550_inst
    process(AND_u1_u1_544_wire, AND_u1_u1_549_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_544_wire, AND_u1_u1_549_wire, tmp_var);
      AND_u1_u1_550_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_449_inst
    process(pkt_priority_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(pkt_priority_buffer, konst_448_wire_constant, tmp_var);
      EQ_u3_u1_449_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_467_inst
    process(pkt_priority_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(pkt_priority_buffer, konst_466_wire_constant, tmp_var);
      EQ_u3_u1_467_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_485_inst
    process(pkt_priority_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(pkt_priority_buffer, konst_484_wire_constant, tmp_var);
      EQ_u3_u1_485_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_503_inst
    process(pkt_priority_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(pkt_priority_buffer, konst_502_wire_constant, tmp_var);
      EQ_u3_u1_503_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_441_inst
    process(down_counter_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(down_counter_buffer, konst_440_wire_constant, tmp_var);
      d0_442 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_451_inst
    process(p4_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_buffer, tmp_var);
      NOT_u1_u1_451_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_453_inst
    process(p2_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_buffer, tmp_var);
      NOT_u1_u1_453_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_456_inst
    process(p3_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_buffer, tmp_var);
      NOT_u1_u1_456_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_469_inst
    process(p4_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_buffer, tmp_var);
      NOT_u1_u1_469_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_471_inst
    process(p1_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_buffer, tmp_var);
      NOT_u1_u1_471_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_474_inst
    process(p3_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_buffer, tmp_var);
      NOT_u1_u1_474_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_487_inst
    process(p4_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_buffer, tmp_var);
      NOT_u1_u1_487_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_489_inst
    process(p2_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_buffer, tmp_var);
      NOT_u1_u1_489_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_492_inst
    process(p1_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_buffer, tmp_var);
      NOT_u1_u1_492_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_505_inst
    process(p1_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_buffer, tmp_var);
      NOT_u1_u1_505_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_507_inst
    process(p2_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_buffer, tmp_var);
      NOT_u1_u1_507_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_510_inst
    process(p3_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_buffer, tmp_var);
      NOT_u1_u1_510_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_517_inst
    process(d0_442) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", d0_442, tmp_var);
      NOT_u1_u1_517_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_541_inst
    process(select_1_460) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", select_1_460, tmp_var);
      NOT_u1_u1_541_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_543_inst
    process(select_2_478) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", select_2_478, tmp_var);
      NOT_u1_u1_543_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_546_inst
    process(select_3_496) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", select_3_496, tmp_var);
      NOT_u1_u1_546_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_548_inst
    process(select_4_514) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", select_4_514, tmp_var);
      NOT_u1_u1_548_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_559_inst
    process(d0_442) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", d0_442, tmp_var);
      NOT_u1_u1_559_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_458_inst
    process(EQ_u3_u1_449_wire, AND_u1_u1_457_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u3_u1_449_wire, AND_u1_u1_457_wire, tmp_var);
      OR_u1_u1_458_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_476_inst
    process(EQ_u3_u1_467_wire, AND_u1_u1_475_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u3_u1_467_wire, AND_u1_u1_475_wire, tmp_var);
      OR_u1_u1_476_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_494_inst
    process(EQ_u3_u1_485_wire, AND_u1_u1_493_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u3_u1_485_wire, AND_u1_u1_493_wire, tmp_var);
      OR_u1_u1_494_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_512_inst
    process(EQ_u3_u1_503_wire, AND_u1_u1_511_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u3_u1_503_wire, AND_u1_u1_511_wire, tmp_var);
      OR_u1_u1_512_wire <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_525_inst
    process(MUX_520_wire, MUX_524_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_520_wire, MUX_524_wire, tmp_var);
      OR_u3_u3_525_wire <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_530_inst
    process(OR_u3_u3_525_wire, MUX_529_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u3_u3_525_wire, MUX_529_wire, tmp_var);
      OR_u3_u3_530_wire <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_539_inst
    process(MUX_534_wire, MUX_538_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_534_wire, MUX_538_wire, tmp_var);
      OR_u3_u3_539_wire <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_554_inst
    process(OR_u3_u3_539_wire, MUX_553_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u3_u3_539_wire, MUX_553_wire, tmp_var);
      OR_u3_u3_554_wire <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_555_inst
    process(OR_u3_u3_530_wire, OR_u3_u3_554_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u3_u3_530_wire, OR_u3_u3_554_wire, tmp_var);
      next_active_packet_buffer <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_567_inst
    process(MUX_562_wire, MUX_566_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_562_wire, MUX_566_wire, tmp_var);
      OR_u3_u3_567_wire <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_572_inst
    process(OR_u3_u3_567_wire, MUX_571_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u3_u3_567_wire, MUX_571_wire, tmp_var);
      OR_u3_u3_572_wire <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_581_inst
    process(MUX_576_wire, MUX_580_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_576_wire, MUX_580_wire, tmp_var);
      OR_u3_u3_581_wire <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_582_inst
    process(OR_u3_u3_572_wire, OR_u3_u3_581_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u3_u3_572_wire, OR_u3_u3_581_wire, tmp_var);
      next_pkt_priority_buffer <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end prioritySelect_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    in_data_1_pipe_write_data: in std_logic_vector(31 downto 0);
    in_data_1_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_1_pipe_write_ack : out std_logic_vector(0 downto 0);
    in_data_2_pipe_write_data: in std_logic_vector(31 downto 0);
    in_data_2_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_2_pipe_write_ack : out std_logic_vector(0 downto 0);
    in_data_3_pipe_write_data: in std_logic_vector(31 downto 0);
    in_data_3_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_3_pipe_write_ack : out std_logic_vector(0 downto 0);
    in_data_4_pipe_write_data: in std_logic_vector(31 downto 0);
    in_data_4_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_4_pipe_write_ack : out std_logic_vector(0 downto 0);
    out_data_1_pipe_read_data: out std_logic_vector(31 downto 0);
    out_data_1_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_1_pipe_read_ack : out std_logic_vector(0 downto 0);
    out_data_2_pipe_read_data: out std_logic_vector(31 downto 0);
    out_data_2_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_2_pipe_read_ack : out std_logic_vector(0 downto 0);
    out_data_3_pipe_read_data: out std_logic_vector(31 downto 0);
    out_data_3_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_3_pipe_read_ack : out std_logic_vector(0 downto 0);
    out_data_4_pipe_read_data: out std_logic_vector(31 downto 0);
    out_data_4_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_4_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- declarations related to module inputPort_1_Daemon
  component inputPort_1_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      in_data_1_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_1_pipe_read_data : in   std_logic_vector(31 downto 0);
      noblock_obuf_1_3_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_3_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_1_4_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_4_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_1_1_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_1_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_1_2_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_2_pipe_write_data : out  std_logic_vector(32 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module inputPort_1_Daemon
  signal inputPort_1_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal inputPort_1_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal inputPort_1_Daemon_start_req : std_logic;
  signal inputPort_1_Daemon_start_ack : std_logic;
  signal inputPort_1_Daemon_fin_req   : std_logic;
  signal inputPort_1_Daemon_fin_ack : std_logic;
  -- declarations related to module inputPort_2_Daemon
  component inputPort_2_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      in_data_2_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_2_pipe_read_data : in   std_logic_vector(31 downto 0);
      noblock_obuf_2_1_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_1_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_2_2_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_2_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_2_3_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_3_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_2_4_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_4_pipe_write_data : out  std_logic_vector(32 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module inputPort_2_Daemon
  signal inputPort_2_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal inputPort_2_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal inputPort_2_Daemon_start_req : std_logic;
  signal inputPort_2_Daemon_start_ack : std_logic;
  signal inputPort_2_Daemon_fin_req   : std_logic;
  signal inputPort_2_Daemon_fin_ack : std_logic;
  -- declarations related to module inputPort_3_Daemon
  component inputPort_3_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      in_data_3_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_3_pipe_read_data : in   std_logic_vector(31 downto 0);
      noblock_obuf_3_2_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_2_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_3_3_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_3_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_3_4_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_4_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_3_1_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_1_pipe_write_data : out  std_logic_vector(32 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module inputPort_3_Daemon
  signal inputPort_3_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal inputPort_3_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal inputPort_3_Daemon_start_req : std_logic;
  signal inputPort_3_Daemon_start_ack : std_logic;
  signal inputPort_3_Daemon_fin_req   : std_logic;
  signal inputPort_3_Daemon_fin_ack : std_logic;
  -- declarations related to module inputPort_4_Daemon
  component inputPort_4_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      in_data_4_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_4_pipe_read_data : in   std_logic_vector(31 downto 0);
      noblock_obuf_4_1_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_1_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_4_2_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_2_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_4_3_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_3_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_4_4_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_4_pipe_write_data : out  std_logic_vector(32 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module inputPort_4_Daemon
  signal inputPort_4_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal inputPort_4_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal inputPort_4_Daemon_start_req : std_logic;
  signal inputPort_4_Daemon_start_ack : std_logic;
  signal inputPort_4_Daemon_fin_req   : std_logic;
  signal inputPort_4_Daemon_fin_ack : std_logic;
  -- declarations related to module outputPort_1_Daemon
  component outputPort_1_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      noblock_obuf_4_1_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_1_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_2_1_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_1_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_1_1_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_1_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_3_1_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_1_pipe_read_data : in   std_logic_vector(32 downto 0);
      out_data_1_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_1_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module outputPort_1_Daemon
  signal outputPort_1_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal outputPort_1_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal outputPort_1_Daemon_start_req : std_logic;
  signal outputPort_1_Daemon_start_ack : std_logic;
  signal outputPort_1_Daemon_fin_req   : std_logic;
  signal outputPort_1_Daemon_fin_ack : std_logic;
  -- declarations related to module outputPort_2_Daemon
  component outputPort_2_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      noblock_obuf_1_2_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_2_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_3_2_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_2_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_4_2_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_2_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_2_2_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_2_pipe_read_data : in   std_logic_vector(32 downto 0);
      out_data_2_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_2_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module outputPort_2_Daemon
  signal outputPort_2_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal outputPort_2_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal outputPort_2_Daemon_start_req : std_logic;
  signal outputPort_2_Daemon_start_ack : std_logic;
  signal outputPort_2_Daemon_fin_req   : std_logic;
  signal outputPort_2_Daemon_fin_ack : std_logic;
  -- declarations related to module outputPort_3_Daemon
  component outputPort_3_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      noblock_obuf_1_3_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_3_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_3_3_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_3_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_4_3_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_3_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_2_3_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_3_pipe_read_data : in   std_logic_vector(32 downto 0);
      out_data_3_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_3_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module outputPort_3_Daemon
  signal outputPort_3_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal outputPort_3_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal outputPort_3_Daemon_start_req : std_logic;
  signal outputPort_3_Daemon_start_ack : std_logic;
  signal outputPort_3_Daemon_fin_req   : std_logic;
  signal outputPort_3_Daemon_fin_ack : std_logic;
  -- declarations related to module outputPort_4_Daemon
  component outputPort_4_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      noblock_obuf_1_4_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_4_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_3_4_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_4_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_2_4_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_4_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_4_4_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_4_pipe_read_data : in   std_logic_vector(32 downto 0);
      out_data_4_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_4_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module outputPort_4_Daemon
  signal outputPort_4_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal outputPort_4_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal outputPort_4_Daemon_start_req : std_logic;
  signal outputPort_4_Daemon_start_ack : std_logic;
  signal outputPort_4_Daemon_fin_req   : std_logic;
  signal outputPort_4_Daemon_fin_ack : std_logic;
  -- declarations related to module prioritySelect
  -- aggregate signals for read from pipe in_data_1
  signal in_data_1_pipe_read_data: std_logic_vector(31 downto 0);
  signal in_data_1_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_data_2
  signal in_data_2_pipe_read_data: std_logic_vector(31 downto 0);
  signal in_data_2_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_data_3
  signal in_data_3_pipe_read_data: std_logic_vector(31 downto 0);
  signal in_data_3_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_data_4
  signal in_data_4_pipe_read_data: std_logic_vector(31 downto 0);
  signal in_data_4_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_4_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_1_1
  signal noblock_obuf_1_1_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_1_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_1_1
  signal noblock_obuf_1_1_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_1_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_1_2
  signal noblock_obuf_1_2_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_2_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_1_2
  signal noblock_obuf_1_2_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_2_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_1_3
  signal noblock_obuf_1_3_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_3_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_1_3
  signal noblock_obuf_1_3_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_3_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_1_4
  signal noblock_obuf_1_4_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_4_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_4_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_1_4
  signal noblock_obuf_1_4_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_4_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_4_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_2_1
  signal noblock_obuf_2_1_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_1_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_2_1
  signal noblock_obuf_2_1_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_1_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_2_2
  signal noblock_obuf_2_2_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_2_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_2_2
  signal noblock_obuf_2_2_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_2_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_2_3
  signal noblock_obuf_2_3_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_3_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_2_3
  signal noblock_obuf_2_3_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_3_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_2_4
  signal noblock_obuf_2_4_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_4_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_4_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_2_4
  signal noblock_obuf_2_4_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_4_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_4_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_3_1
  signal noblock_obuf_3_1_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_1_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_3_1
  signal noblock_obuf_3_1_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_1_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_3_2
  signal noblock_obuf_3_2_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_2_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_3_2
  signal noblock_obuf_3_2_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_2_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_3_3
  signal noblock_obuf_3_3_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_3_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_3_3
  signal noblock_obuf_3_3_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_3_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_3_4
  signal noblock_obuf_3_4_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_4_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_4_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_3_4
  signal noblock_obuf_3_4_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_4_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_4_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_4_1
  signal noblock_obuf_4_1_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_1_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_4_1
  signal noblock_obuf_4_1_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_1_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_4_2
  signal noblock_obuf_4_2_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_2_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_4_2
  signal noblock_obuf_4_2_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_2_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_4_3
  signal noblock_obuf_4_3_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_3_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_4_3
  signal noblock_obuf_4_3_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_3_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_4_4
  signal noblock_obuf_4_4_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_4_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_4_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_4_4
  signal noblock_obuf_4_4_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_4_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_4_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data_1
  signal out_data_1_pipe_write_data: std_logic_vector(31 downto 0);
  signal out_data_1_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data_2
  signal out_data_2_pipe_write_data: std_logic_vector(31 downto 0);
  signal out_data_2_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data_3
  signal out_data_3_pipe_write_data: std_logic_vector(31 downto 0);
  signal out_data_3_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data_4
  signal out_data_4_pipe_write_data: std_logic_vector(31 downto 0);
  signal out_data_4_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_4_pipe_write_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module inputPort_1_Daemon
  inputPort_1_Daemon_instance:inputPort_1_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => inputPort_1_Daemon_start_req,
      start_ack => inputPort_1_Daemon_start_ack,
      fin_req => inputPort_1_Daemon_fin_req,
      fin_ack => inputPort_1_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      in_data_1_pipe_read_req => in_data_1_pipe_read_req(0 downto 0),
      in_data_1_pipe_read_ack => in_data_1_pipe_read_ack(0 downto 0),
      in_data_1_pipe_read_data => in_data_1_pipe_read_data(31 downto 0),
      noblock_obuf_1_3_pipe_write_req => noblock_obuf_1_3_pipe_write_req(0 downto 0),
      noblock_obuf_1_3_pipe_write_ack => noblock_obuf_1_3_pipe_write_ack(0 downto 0),
      noblock_obuf_1_3_pipe_write_data => noblock_obuf_1_3_pipe_write_data(32 downto 0),
      noblock_obuf_1_4_pipe_write_req => noblock_obuf_1_4_pipe_write_req(0 downto 0),
      noblock_obuf_1_4_pipe_write_ack => noblock_obuf_1_4_pipe_write_ack(0 downto 0),
      noblock_obuf_1_4_pipe_write_data => noblock_obuf_1_4_pipe_write_data(32 downto 0),
      noblock_obuf_1_1_pipe_write_req => noblock_obuf_1_1_pipe_write_req(0 downto 0),
      noblock_obuf_1_1_pipe_write_ack => noblock_obuf_1_1_pipe_write_ack(0 downto 0),
      noblock_obuf_1_1_pipe_write_data => noblock_obuf_1_1_pipe_write_data(32 downto 0),
      noblock_obuf_1_2_pipe_write_req => noblock_obuf_1_2_pipe_write_req(0 downto 0),
      noblock_obuf_1_2_pipe_write_ack => noblock_obuf_1_2_pipe_write_ack(0 downto 0),
      noblock_obuf_1_2_pipe_write_data => noblock_obuf_1_2_pipe_write_data(32 downto 0),
      tag_in => inputPort_1_Daemon_tag_in,
      tag_out => inputPort_1_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  inputPort_1_Daemon_tag_in <= (others => '0');
  inputPort_1_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => inputPort_1_Daemon_start_req, start_ack => inputPort_1_Daemon_start_ack,  fin_req => inputPort_1_Daemon_fin_req,  fin_ack => inputPort_1_Daemon_fin_ack);
  -- module inputPort_2_Daemon
  inputPort_2_Daemon_instance:inputPort_2_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => inputPort_2_Daemon_start_req,
      start_ack => inputPort_2_Daemon_start_ack,
      fin_req => inputPort_2_Daemon_fin_req,
      fin_ack => inputPort_2_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      in_data_2_pipe_read_req => in_data_2_pipe_read_req(0 downto 0),
      in_data_2_pipe_read_ack => in_data_2_pipe_read_ack(0 downto 0),
      in_data_2_pipe_read_data => in_data_2_pipe_read_data(31 downto 0),
      noblock_obuf_2_1_pipe_write_req => noblock_obuf_2_1_pipe_write_req(0 downto 0),
      noblock_obuf_2_1_pipe_write_ack => noblock_obuf_2_1_pipe_write_ack(0 downto 0),
      noblock_obuf_2_1_pipe_write_data => noblock_obuf_2_1_pipe_write_data(32 downto 0),
      noblock_obuf_2_2_pipe_write_req => noblock_obuf_2_2_pipe_write_req(0 downto 0),
      noblock_obuf_2_2_pipe_write_ack => noblock_obuf_2_2_pipe_write_ack(0 downto 0),
      noblock_obuf_2_2_pipe_write_data => noblock_obuf_2_2_pipe_write_data(32 downto 0),
      noblock_obuf_2_3_pipe_write_req => noblock_obuf_2_3_pipe_write_req(0 downto 0),
      noblock_obuf_2_3_pipe_write_ack => noblock_obuf_2_3_pipe_write_ack(0 downto 0),
      noblock_obuf_2_3_pipe_write_data => noblock_obuf_2_3_pipe_write_data(32 downto 0),
      noblock_obuf_2_4_pipe_write_req => noblock_obuf_2_4_pipe_write_req(0 downto 0),
      noblock_obuf_2_4_pipe_write_ack => noblock_obuf_2_4_pipe_write_ack(0 downto 0),
      noblock_obuf_2_4_pipe_write_data => noblock_obuf_2_4_pipe_write_data(32 downto 0),
      tag_in => inputPort_2_Daemon_tag_in,
      tag_out => inputPort_2_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  inputPort_2_Daemon_tag_in <= (others => '0');
  inputPort_2_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => inputPort_2_Daemon_start_req, start_ack => inputPort_2_Daemon_start_ack,  fin_req => inputPort_2_Daemon_fin_req,  fin_ack => inputPort_2_Daemon_fin_ack);
  -- module inputPort_3_Daemon
  inputPort_3_Daemon_instance:inputPort_3_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => inputPort_3_Daemon_start_req,
      start_ack => inputPort_3_Daemon_start_ack,
      fin_req => inputPort_3_Daemon_fin_req,
      fin_ack => inputPort_3_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      in_data_3_pipe_read_req => in_data_3_pipe_read_req(0 downto 0),
      in_data_3_pipe_read_ack => in_data_3_pipe_read_ack(0 downto 0),
      in_data_3_pipe_read_data => in_data_3_pipe_read_data(31 downto 0),
      noblock_obuf_3_2_pipe_write_req => noblock_obuf_3_2_pipe_write_req(0 downto 0),
      noblock_obuf_3_2_pipe_write_ack => noblock_obuf_3_2_pipe_write_ack(0 downto 0),
      noblock_obuf_3_2_pipe_write_data => noblock_obuf_3_2_pipe_write_data(32 downto 0),
      noblock_obuf_3_3_pipe_write_req => noblock_obuf_3_3_pipe_write_req(0 downto 0),
      noblock_obuf_3_3_pipe_write_ack => noblock_obuf_3_3_pipe_write_ack(0 downto 0),
      noblock_obuf_3_3_pipe_write_data => noblock_obuf_3_3_pipe_write_data(32 downto 0),
      noblock_obuf_3_4_pipe_write_req => noblock_obuf_3_4_pipe_write_req(0 downto 0),
      noblock_obuf_3_4_pipe_write_ack => noblock_obuf_3_4_pipe_write_ack(0 downto 0),
      noblock_obuf_3_4_pipe_write_data => noblock_obuf_3_4_pipe_write_data(32 downto 0),
      noblock_obuf_3_1_pipe_write_req => noblock_obuf_3_1_pipe_write_req(0 downto 0),
      noblock_obuf_3_1_pipe_write_ack => noblock_obuf_3_1_pipe_write_ack(0 downto 0),
      noblock_obuf_3_1_pipe_write_data => noblock_obuf_3_1_pipe_write_data(32 downto 0),
      tag_in => inputPort_3_Daemon_tag_in,
      tag_out => inputPort_3_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  inputPort_3_Daemon_tag_in <= (others => '0');
  inputPort_3_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => inputPort_3_Daemon_start_req, start_ack => inputPort_3_Daemon_start_ack,  fin_req => inputPort_3_Daemon_fin_req,  fin_ack => inputPort_3_Daemon_fin_ack);
  -- module inputPort_4_Daemon
  inputPort_4_Daemon_instance:inputPort_4_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => inputPort_4_Daemon_start_req,
      start_ack => inputPort_4_Daemon_start_ack,
      fin_req => inputPort_4_Daemon_fin_req,
      fin_ack => inputPort_4_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      in_data_4_pipe_read_req => in_data_4_pipe_read_req(0 downto 0),
      in_data_4_pipe_read_ack => in_data_4_pipe_read_ack(0 downto 0),
      in_data_4_pipe_read_data => in_data_4_pipe_read_data(31 downto 0),
      noblock_obuf_4_1_pipe_write_req => noblock_obuf_4_1_pipe_write_req(0 downto 0),
      noblock_obuf_4_1_pipe_write_ack => noblock_obuf_4_1_pipe_write_ack(0 downto 0),
      noblock_obuf_4_1_pipe_write_data => noblock_obuf_4_1_pipe_write_data(32 downto 0),
      noblock_obuf_4_2_pipe_write_req => noblock_obuf_4_2_pipe_write_req(0 downto 0),
      noblock_obuf_4_2_pipe_write_ack => noblock_obuf_4_2_pipe_write_ack(0 downto 0),
      noblock_obuf_4_2_pipe_write_data => noblock_obuf_4_2_pipe_write_data(32 downto 0),
      noblock_obuf_4_3_pipe_write_req => noblock_obuf_4_3_pipe_write_req(0 downto 0),
      noblock_obuf_4_3_pipe_write_ack => noblock_obuf_4_3_pipe_write_ack(0 downto 0),
      noblock_obuf_4_3_pipe_write_data => noblock_obuf_4_3_pipe_write_data(32 downto 0),
      noblock_obuf_4_4_pipe_write_req => noblock_obuf_4_4_pipe_write_req(0 downto 0),
      noblock_obuf_4_4_pipe_write_ack => noblock_obuf_4_4_pipe_write_ack(0 downto 0),
      noblock_obuf_4_4_pipe_write_data => noblock_obuf_4_4_pipe_write_data(32 downto 0),
      tag_in => inputPort_4_Daemon_tag_in,
      tag_out => inputPort_4_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  inputPort_4_Daemon_tag_in <= (others => '0');
  inputPort_4_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => inputPort_4_Daemon_start_req, start_ack => inputPort_4_Daemon_start_ack,  fin_req => inputPort_4_Daemon_fin_req,  fin_ack => inputPort_4_Daemon_fin_ack);
  -- module outputPort_1_Daemon
  outputPort_1_Daemon_instance:outputPort_1_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => outputPort_1_Daemon_start_req,
      start_ack => outputPort_1_Daemon_start_ack,
      fin_req => outputPort_1_Daemon_fin_req,
      fin_ack => outputPort_1_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      noblock_obuf_4_1_pipe_read_req => noblock_obuf_4_1_pipe_read_req(0 downto 0),
      noblock_obuf_4_1_pipe_read_ack => noblock_obuf_4_1_pipe_read_ack(0 downto 0),
      noblock_obuf_4_1_pipe_read_data => noblock_obuf_4_1_pipe_read_data(32 downto 0),
      noblock_obuf_2_1_pipe_read_req => noblock_obuf_2_1_pipe_read_req(0 downto 0),
      noblock_obuf_2_1_pipe_read_ack => noblock_obuf_2_1_pipe_read_ack(0 downto 0),
      noblock_obuf_2_1_pipe_read_data => noblock_obuf_2_1_pipe_read_data(32 downto 0),
      noblock_obuf_1_1_pipe_read_req => noblock_obuf_1_1_pipe_read_req(0 downto 0),
      noblock_obuf_1_1_pipe_read_ack => noblock_obuf_1_1_pipe_read_ack(0 downto 0),
      noblock_obuf_1_1_pipe_read_data => noblock_obuf_1_1_pipe_read_data(32 downto 0),
      noblock_obuf_3_1_pipe_read_req => noblock_obuf_3_1_pipe_read_req(0 downto 0),
      noblock_obuf_3_1_pipe_read_ack => noblock_obuf_3_1_pipe_read_ack(0 downto 0),
      noblock_obuf_3_1_pipe_read_data => noblock_obuf_3_1_pipe_read_data(32 downto 0),
      out_data_1_pipe_write_req => out_data_1_pipe_write_req(0 downto 0),
      out_data_1_pipe_write_ack => out_data_1_pipe_write_ack(0 downto 0),
      out_data_1_pipe_write_data => out_data_1_pipe_write_data(31 downto 0),
      tag_in => outputPort_1_Daemon_tag_in,
      tag_out => outputPort_1_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  outputPort_1_Daemon_tag_in <= (others => '0');
  outputPort_1_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => outputPort_1_Daemon_start_req, start_ack => outputPort_1_Daemon_start_ack,  fin_req => outputPort_1_Daemon_fin_req,  fin_ack => outputPort_1_Daemon_fin_ack);
  -- module outputPort_2_Daemon
  outputPort_2_Daemon_instance:outputPort_2_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => outputPort_2_Daemon_start_req,
      start_ack => outputPort_2_Daemon_start_ack,
      fin_req => outputPort_2_Daemon_fin_req,
      fin_ack => outputPort_2_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      noblock_obuf_1_2_pipe_read_req => noblock_obuf_1_2_pipe_read_req(0 downto 0),
      noblock_obuf_1_2_pipe_read_ack => noblock_obuf_1_2_pipe_read_ack(0 downto 0),
      noblock_obuf_1_2_pipe_read_data => noblock_obuf_1_2_pipe_read_data(32 downto 0),
      noblock_obuf_3_2_pipe_read_req => noblock_obuf_3_2_pipe_read_req(0 downto 0),
      noblock_obuf_3_2_pipe_read_ack => noblock_obuf_3_2_pipe_read_ack(0 downto 0),
      noblock_obuf_3_2_pipe_read_data => noblock_obuf_3_2_pipe_read_data(32 downto 0),
      noblock_obuf_4_2_pipe_read_req => noblock_obuf_4_2_pipe_read_req(0 downto 0),
      noblock_obuf_4_2_pipe_read_ack => noblock_obuf_4_2_pipe_read_ack(0 downto 0),
      noblock_obuf_4_2_pipe_read_data => noblock_obuf_4_2_pipe_read_data(32 downto 0),
      noblock_obuf_2_2_pipe_read_req => noblock_obuf_2_2_pipe_read_req(0 downto 0),
      noblock_obuf_2_2_pipe_read_ack => noblock_obuf_2_2_pipe_read_ack(0 downto 0),
      noblock_obuf_2_2_pipe_read_data => noblock_obuf_2_2_pipe_read_data(32 downto 0),
      out_data_2_pipe_write_req => out_data_2_pipe_write_req(0 downto 0),
      out_data_2_pipe_write_ack => out_data_2_pipe_write_ack(0 downto 0),
      out_data_2_pipe_write_data => out_data_2_pipe_write_data(31 downto 0),
      tag_in => outputPort_2_Daemon_tag_in,
      tag_out => outputPort_2_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  outputPort_2_Daemon_tag_in <= (others => '0');
  outputPort_2_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => outputPort_2_Daemon_start_req, start_ack => outputPort_2_Daemon_start_ack,  fin_req => outputPort_2_Daemon_fin_req,  fin_ack => outputPort_2_Daemon_fin_ack);
  -- module outputPort_3_Daemon
  outputPort_3_Daemon_instance:outputPort_3_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => outputPort_3_Daemon_start_req,
      start_ack => outputPort_3_Daemon_start_ack,
      fin_req => outputPort_3_Daemon_fin_req,
      fin_ack => outputPort_3_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      noblock_obuf_1_3_pipe_read_req => noblock_obuf_1_3_pipe_read_req(0 downto 0),
      noblock_obuf_1_3_pipe_read_ack => noblock_obuf_1_3_pipe_read_ack(0 downto 0),
      noblock_obuf_1_3_pipe_read_data => noblock_obuf_1_3_pipe_read_data(32 downto 0),
      noblock_obuf_3_3_pipe_read_req => noblock_obuf_3_3_pipe_read_req(0 downto 0),
      noblock_obuf_3_3_pipe_read_ack => noblock_obuf_3_3_pipe_read_ack(0 downto 0),
      noblock_obuf_3_3_pipe_read_data => noblock_obuf_3_3_pipe_read_data(32 downto 0),
      noblock_obuf_4_3_pipe_read_req => noblock_obuf_4_3_pipe_read_req(0 downto 0),
      noblock_obuf_4_3_pipe_read_ack => noblock_obuf_4_3_pipe_read_ack(0 downto 0),
      noblock_obuf_4_3_pipe_read_data => noblock_obuf_4_3_pipe_read_data(32 downto 0),
      noblock_obuf_2_3_pipe_read_req => noblock_obuf_2_3_pipe_read_req(0 downto 0),
      noblock_obuf_2_3_pipe_read_ack => noblock_obuf_2_3_pipe_read_ack(0 downto 0),
      noblock_obuf_2_3_pipe_read_data => noblock_obuf_2_3_pipe_read_data(32 downto 0),
      out_data_3_pipe_write_req => out_data_3_pipe_write_req(0 downto 0),
      out_data_3_pipe_write_ack => out_data_3_pipe_write_ack(0 downto 0),
      out_data_3_pipe_write_data => out_data_3_pipe_write_data(31 downto 0),
      tag_in => outputPort_3_Daemon_tag_in,
      tag_out => outputPort_3_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  outputPort_3_Daemon_tag_in <= (others => '0');
  outputPort_3_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => outputPort_3_Daemon_start_req, start_ack => outputPort_3_Daemon_start_ack,  fin_req => outputPort_3_Daemon_fin_req,  fin_ack => outputPort_3_Daemon_fin_ack);
  -- module outputPort_4_Daemon
  outputPort_4_Daemon_instance:outputPort_4_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => outputPort_4_Daemon_start_req,
      start_ack => outputPort_4_Daemon_start_ack,
      fin_req => outputPort_4_Daemon_fin_req,
      fin_ack => outputPort_4_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      noblock_obuf_1_4_pipe_read_req => noblock_obuf_1_4_pipe_read_req(0 downto 0),
      noblock_obuf_1_4_pipe_read_ack => noblock_obuf_1_4_pipe_read_ack(0 downto 0),
      noblock_obuf_1_4_pipe_read_data => noblock_obuf_1_4_pipe_read_data(32 downto 0),
      noblock_obuf_3_4_pipe_read_req => noblock_obuf_3_4_pipe_read_req(0 downto 0),
      noblock_obuf_3_4_pipe_read_ack => noblock_obuf_3_4_pipe_read_ack(0 downto 0),
      noblock_obuf_3_4_pipe_read_data => noblock_obuf_3_4_pipe_read_data(32 downto 0),
      noblock_obuf_2_4_pipe_read_req => noblock_obuf_2_4_pipe_read_req(0 downto 0),
      noblock_obuf_2_4_pipe_read_ack => noblock_obuf_2_4_pipe_read_ack(0 downto 0),
      noblock_obuf_2_4_pipe_read_data => noblock_obuf_2_4_pipe_read_data(32 downto 0),
      noblock_obuf_4_4_pipe_read_req => noblock_obuf_4_4_pipe_read_req(0 downto 0),
      noblock_obuf_4_4_pipe_read_ack => noblock_obuf_4_4_pipe_read_ack(0 downto 0),
      noblock_obuf_4_4_pipe_read_data => noblock_obuf_4_4_pipe_read_data(32 downto 0),
      out_data_4_pipe_write_req => out_data_4_pipe_write_req(0 downto 0),
      out_data_4_pipe_write_ack => out_data_4_pipe_write_ack(0 downto 0),
      out_data_4_pipe_write_data => out_data_4_pipe_write_data(31 downto 0),
      tag_in => outputPort_4_Daemon_tag_in,
      tag_out => outputPort_4_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  outputPort_4_Daemon_tag_in <= (others => '0');
  outputPort_4_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => outputPort_4_Daemon_start_req, start_ack => outputPort_4_Daemon_start_ack,  fin_req => outputPort_4_Daemon_fin_req,  fin_ack => outputPort_4_Daemon_fin_ack);
  in_data_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe in_data_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => in_data_1_pipe_read_req,
      read_ack => in_data_1_pipe_read_ack,
      read_data => in_data_1_pipe_read_data,
      write_req => in_data_1_pipe_write_req,
      write_ack => in_data_1_pipe_write_ack,
      write_data => in_data_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  in_data_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe in_data_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => in_data_2_pipe_read_req,
      read_ack => in_data_2_pipe_read_ack,
      read_data => in_data_2_pipe_read_data,
      write_req => in_data_2_pipe_write_req,
      write_ack => in_data_2_pipe_write_ack,
      write_data => in_data_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  in_data_3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe in_data_3",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => in_data_3_pipe_read_req,
      read_ack => in_data_3_pipe_read_ack,
      read_data => in_data_3_pipe_read_data,
      write_req => in_data_3_pipe_write_req,
      write_ack => in_data_3_pipe_write_ack,
      write_data => in_data_3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  in_data_4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe in_data_4",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => in_data_4_pipe_read_req,
      read_ack => in_data_4_pipe_read_ack,
      read_data => in_data_4_pipe_read_data,
      write_req => in_data_4_pipe_write_req,
      write_ack => in_data_4_pipe_write_ack,
      write_data => in_data_4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_1_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_1_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_1_1_pipe_read_req,
      read_ack => noblock_obuf_1_1_pipe_read_ack,
      read_data => noblock_obuf_1_1_pipe_read_data,
      write_req => noblock_obuf_1_1_pipe_write_req,
      write_ack => noblock_obuf_1_1_pipe_write_ack,
      write_data => noblock_obuf_1_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_1_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_1_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_1_2_pipe_read_req,
      read_ack => noblock_obuf_1_2_pipe_read_ack,
      read_data => noblock_obuf_1_2_pipe_read_data,
      write_req => noblock_obuf_1_2_pipe_write_req,
      write_ack => noblock_obuf_1_2_pipe_write_ack,
      write_data => noblock_obuf_1_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_1_3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_1_3",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_1_3_pipe_read_req,
      read_ack => noblock_obuf_1_3_pipe_read_ack,
      read_data => noblock_obuf_1_3_pipe_read_data,
      write_req => noblock_obuf_1_3_pipe_write_req,
      write_ack => noblock_obuf_1_3_pipe_write_ack,
      write_data => noblock_obuf_1_3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_1_4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_1_4",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_1_4_pipe_read_req,
      read_ack => noblock_obuf_1_4_pipe_read_ack,
      read_data => noblock_obuf_1_4_pipe_read_data,
      write_req => noblock_obuf_1_4_pipe_write_req,
      write_ack => noblock_obuf_1_4_pipe_write_ack,
      write_data => noblock_obuf_1_4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_2_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_2_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_2_1_pipe_read_req,
      read_ack => noblock_obuf_2_1_pipe_read_ack,
      read_data => noblock_obuf_2_1_pipe_read_data,
      write_req => noblock_obuf_2_1_pipe_write_req,
      write_ack => noblock_obuf_2_1_pipe_write_ack,
      write_data => noblock_obuf_2_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_2_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_2_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_2_2_pipe_read_req,
      read_ack => noblock_obuf_2_2_pipe_read_ack,
      read_data => noblock_obuf_2_2_pipe_read_data,
      write_req => noblock_obuf_2_2_pipe_write_req,
      write_ack => noblock_obuf_2_2_pipe_write_ack,
      write_data => noblock_obuf_2_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_2_3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_2_3",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_2_3_pipe_read_req,
      read_ack => noblock_obuf_2_3_pipe_read_ack,
      read_data => noblock_obuf_2_3_pipe_read_data,
      write_req => noblock_obuf_2_3_pipe_write_req,
      write_ack => noblock_obuf_2_3_pipe_write_ack,
      write_data => noblock_obuf_2_3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_2_4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_2_4",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_2_4_pipe_read_req,
      read_ack => noblock_obuf_2_4_pipe_read_ack,
      read_data => noblock_obuf_2_4_pipe_read_data,
      write_req => noblock_obuf_2_4_pipe_write_req,
      write_ack => noblock_obuf_2_4_pipe_write_ack,
      write_data => noblock_obuf_2_4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_3_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_3_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_3_1_pipe_read_req,
      read_ack => noblock_obuf_3_1_pipe_read_ack,
      read_data => noblock_obuf_3_1_pipe_read_data,
      write_req => noblock_obuf_3_1_pipe_write_req,
      write_ack => noblock_obuf_3_1_pipe_write_ack,
      write_data => noblock_obuf_3_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_3_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_3_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_3_2_pipe_read_req,
      read_ack => noblock_obuf_3_2_pipe_read_ack,
      read_data => noblock_obuf_3_2_pipe_read_data,
      write_req => noblock_obuf_3_2_pipe_write_req,
      write_ack => noblock_obuf_3_2_pipe_write_ack,
      write_data => noblock_obuf_3_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_3_3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_3_3",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_3_3_pipe_read_req,
      read_ack => noblock_obuf_3_3_pipe_read_ack,
      read_data => noblock_obuf_3_3_pipe_read_data,
      write_req => noblock_obuf_3_3_pipe_write_req,
      write_ack => noblock_obuf_3_3_pipe_write_ack,
      write_data => noblock_obuf_3_3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_3_4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_3_4",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_3_4_pipe_read_req,
      read_ack => noblock_obuf_3_4_pipe_read_ack,
      read_data => noblock_obuf_3_4_pipe_read_data,
      write_req => noblock_obuf_3_4_pipe_write_req,
      write_ack => noblock_obuf_3_4_pipe_write_ack,
      write_data => noblock_obuf_3_4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_4_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_4_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_4_1_pipe_read_req,
      read_ack => noblock_obuf_4_1_pipe_read_ack,
      read_data => noblock_obuf_4_1_pipe_read_data,
      write_req => noblock_obuf_4_1_pipe_write_req,
      write_ack => noblock_obuf_4_1_pipe_write_ack,
      write_data => noblock_obuf_4_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_4_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_4_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_4_2_pipe_read_req,
      read_ack => noblock_obuf_4_2_pipe_read_ack,
      read_data => noblock_obuf_4_2_pipe_read_data,
      write_req => noblock_obuf_4_2_pipe_write_req,
      write_ack => noblock_obuf_4_2_pipe_write_ack,
      write_data => noblock_obuf_4_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_4_3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_4_3",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_4_3_pipe_read_req,
      read_ack => noblock_obuf_4_3_pipe_read_ack,
      read_data => noblock_obuf_4_3_pipe_read_data,
      write_req => noblock_obuf_4_3_pipe_write_req,
      write_ack => noblock_obuf_4_3_pipe_write_ack,
      write_data => noblock_obuf_4_3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_4_4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_4_4",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_4_4_pipe_read_req,
      read_ack => noblock_obuf_4_4_pipe_read_ack,
      read_data => noblock_obuf_4_4_pipe_read_data,
      write_req => noblock_obuf_4_4_pipe_write_req,
      write_ack => noblock_obuf_4_4_pipe_write_ack,
      write_data => noblock_obuf_4_4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe out_data_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => out_data_1_pipe_read_req,
      read_ack => out_data_1_pipe_read_ack,
      read_data => out_data_1_pipe_read_data,
      write_req => out_data_1_pipe_write_req,
      write_ack => out_data_1_pipe_write_ack,
      write_data => out_data_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe out_data_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => out_data_2_pipe_read_req,
      read_ack => out_data_2_pipe_read_ack,
      read_data => out_data_2_pipe_read_data,
      write_req => out_data_2_pipe_write_req,
      write_ack => out_data_2_pipe_write_ack,
      write_data => out_data_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe out_data_3",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => out_data_3_pipe_read_req,
      read_ack => out_data_3_pipe_read_ack,
      read_data => out_data_3_pipe_read_data,
      write_req => out_data_3_pipe_write_req,
      write_ack => out_data_3_pipe_write_ack,
      write_data => out_data_3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe out_data_4",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => out_data_4_pipe_read_req,
      read_ack => out_data_4_pipe_read_ack,
      read_data => out_data_4_pipe_read_data,
      write_req => out_data_4_pipe_write_req,
      write_ack => out_data_4_pipe_write_ack,
      write_data => out_data_4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- 
end ahir_system_arch;
