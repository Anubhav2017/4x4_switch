-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity inputPort_1_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    in_data_1_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_1_pipe_read_data : in   std_logic_vector(31 downto 0);
    noblock_obuf_1_3_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_3_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_1_4_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_4_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_1_1_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_1_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_1_2_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_2_pipe_write_data : out  std_logic_vector(32 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity inputPort_1_Daemon;
architecture inputPort_1_Daemon_arch of inputPort_1_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal inputPort_1_Daemon_CP_3_start: Boolean;
  signal inputPort_1_Daemon_CP_3_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal phi_stmt_67_req_0 : boolean;
  signal do_while_stmt_65_branch_req_0 : boolean;
  signal phi_stmt_76_req_0 : boolean;
  signal phi_stmt_76_ack_0 : boolean;
  signal phi_stmt_67_req_1 : boolean;
  signal phi_stmt_67_ack_0 : boolean;
  signal next_count_down_103_69_buf_req_0 : boolean;
  signal next_count_down_103_69_buf_ack_0 : boolean;
  signal next_count_down_103_69_buf_req_1 : boolean;
  signal next_count_down_103_69_buf_ack_1 : boolean;
  signal RPIPE_in_data_1_75_inst_req_0 : boolean;
  signal RPIPE_in_data_1_75_inst_ack_0 : boolean;
  signal RPIPE_in_data_1_75_inst_req_1 : boolean;
  signal RPIPE_in_data_1_75_inst_ack_1 : boolean;
  signal phi_stmt_76_req_1 : boolean;
  signal next_last_dest_id_109_79_buf_req_0 : boolean;
  signal next_last_dest_id_109_79_buf_ack_0 : boolean;
  signal next_last_dest_id_109_79_buf_req_1 : boolean;
  signal next_last_dest_id_109_79_buf_ack_1 : boolean;
  signal WPIPE_noblock_obuf_1_1_121_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_1_1_121_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_1_1_121_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_1_1_121_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_1_2_130_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_1_2_130_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_1_2_130_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_1_2_130_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_1_3_139_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_1_3_139_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_1_3_139_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_1_3_139_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_1_4_148_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_1_4_148_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_1_4_148_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_1_4_148_inst_ack_1 : boolean;
  signal do_while_stmt_65_branch_ack_0 : boolean;
  signal do_while_stmt_65_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "inputPort_1_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  inputPort_1_Daemon_CP_3_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "inputPort_1_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_1_Daemon_CP_3_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= inputPort_1_Daemon_CP_3_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_1_Daemon_CP_3_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  inputPort_1_Daemon_CP_3: Block -- control-path 
    signal inputPort_1_Daemon_CP_3_elements: BooleanArray(72 downto 0);
    -- 
  begin -- 
    inputPort_1_Daemon_CP_3_elements(0) <= inputPort_1_Daemon_CP_3_start;
    inputPort_1_Daemon_CP_3_symbol <= inputPort_1_Daemon_CP_3_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_64/$entry
      -- CP-element group 0: 	 branch_block_stmt_64/branch_block_stmt_64__entry__
      -- CP-element group 0: 	 branch_block_stmt_64/do_while_stmt_65__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	72 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_64/$exit
      -- CP-element group 1: 	 branch_block_stmt_64/branch_block_stmt_64__exit__
      -- CP-element group 1: 	 branch_block_stmt_64/do_while_stmt_65__exit__
      -- 
    inputPort_1_Daemon_CP_3_elements(1) <= inputPort_1_Daemon_CP_3_elements(72);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_64/do_while_stmt_65/$entry
      -- CP-element group 2: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65__entry__
      -- 
    inputPort_1_Daemon_CP_3_elements(2) <= inputPort_1_Daemon_CP_3_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	72 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65__exit__
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_64/do_while_stmt_65/loop_back
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	70 
    -- CP-element group 5: 	71 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_64/do_while_stmt_65/condition_done
      -- CP-element group 5: 	 branch_block_stmt_64/do_while_stmt_65/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_64/do_while_stmt_65/loop_taken/$entry
      -- 
    inputPort_1_Daemon_CP_3_elements(5) <= inputPort_1_Daemon_CP_3_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	69 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_64/do_while_stmt_65/loop_body_done
      -- 
    inputPort_1_Daemon_CP_3_elements(6) <= inputPort_1_Daemon_CP_3_elements(69);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	43 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/back_edge_to_loop_body
      -- 
    inputPort_1_Daemon_CP_3_elements(7) <= inputPort_1_Daemon_CP_3_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	45 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/first_time_through_loop_body
      -- 
    inputPort_1_Daemon_CP_3_elements(8) <= inputPort_1_Daemon_CP_3_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	37 
    -- CP-element group 9: 	38 
    -- CP-element group 9: 	68 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_73_sample_start_
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	68 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/condition_evaluated
      -- 
    condition_evaluated_27_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_27_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(10), ack => do_while_stmt_65_branch_req_0); -- 
    inputPort_1_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(14) & inputPort_1_Daemon_CP_3_elements(68);
      gj_inputPort_1_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	37 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11: 	39 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_sample_start__ps
      -- 
    inputPort_1_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(9) & inputPort_1_Daemon_CP_3_elements(15) & inputPort_1_Daemon_CP_3_elements(37) & inputPort_1_Daemon_CP_3_elements(14);
      gj_inputPort_1_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	40 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	69 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	37 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_73_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_sample_completed_
      -- 
    inputPort_1_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(17) & inputPort_1_Daemon_CP_3_elements(35) & inputPort_1_Daemon_CP_3_elements(40);
      gj_inputPort_1_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	32 
    -- CP-element group 13: 	38 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13: 	41 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_update_start__ps
      -- 
    inputPort_1_Daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(16) & inputPort_1_Daemon_CP_3_elements(32) & inputPort_1_Daemon_CP_3_elements(38);
      gj_inputPort_1_Daemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	36 
    -- CP-element group 14: 	42 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/aggregated_phi_update_ack
      -- 
    inputPort_1_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(18) & inputPort_1_Daemon_CP_3_elements(36) & inputPort_1_Daemon_CP_3_elements(42);
      gj_inputPort_1_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_sample_start_
      -- 
    inputPort_1_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(9) & inputPort_1_Daemon_CP_3_elements(12);
      gj_inputPort_1_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	57 
    -- CP-element group 16: 	60 
    -- CP-element group 16: 	63 
    -- CP-element group 16: 	66 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_update_start_
      -- 
    inputPort_1_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(9) & inputPort_1_Daemon_CP_3_elements(57) & inputPort_1_Daemon_CP_3_elements(60) & inputPort_1_Daemon_CP_3_elements(63) & inputPort_1_Daemon_CP_3_elements(66);
      gj_inputPort_1_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_sample_completed__ps
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	56 
    -- CP-element group 18: 	59 
    -- CP-element group 18: 	62 
    -- CP-element group 18: 	65 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_update_completed__ps
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_loopback_trigger
      -- 
    inputPort_1_Daemon_CP_3_elements(19) <= inputPort_1_Daemon_CP_3_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_loopback_sample_req_ps
      -- 
    phi_stmt_67_loopback_sample_req_42_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_67_loopback_sample_req_42_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(20), ack => phi_stmt_67_req_0); -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_entry_trigger
      -- 
    inputPort_1_Daemon_CP_3_elements(21) <= inputPort_1_Daemon_CP_3_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_entry_sample_req_ps
      -- 
    phi_stmt_67_entry_sample_req_45_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_67_entry_sample_req_45_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(22), ack => phi_stmt_67_req_1); -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_67_phi_mux_ack_ps
      -- 
    phi_stmt_67_phi_mux_ack_48_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_67_ack_0, ack => inputPort_1_Daemon_CP_3_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_69_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_69_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_69_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_69_Sample/req
      -- 
    req_61_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_61_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(24), ack => next_count_down_103_69_buf_req_0); -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_69_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_69_update_start_
      -- CP-element group 25: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_69_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_69_Update/req
      -- 
    req_66_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_66_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(25), ack => next_count_down_103_69_buf_req_1); -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_69_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_69_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_69_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_69_Sample/ack
      -- 
    ack_62_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_103_69_buf_ack_0, ack => inputPort_1_Daemon_CP_3_elements(26)); -- 
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_69_update_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_69_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_69_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_count_down_69_Update/ack
      -- 
    ack_67_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_103_69_buf_ack_1, ack => inputPort_1_Daemon_CP_3_elements(27)); -- 
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/type_cast_72_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/type_cast_72_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/type_cast_72_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/type_cast_72_sample_completed_
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/type_cast_72_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/type_cast_72_update_start_
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/type_cast_72_update_completed__ps
      -- 
    inputPort_1_Daemon_CP_3_elements(30) <= inputPort_1_Daemon_CP_3_elements(31);
    -- CP-element group 31:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	30 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/type_cast_72_update_completed_
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(31) is a control-delay.
    cp_element_31_delay: control_delay_element  generic map(name => " 31_delay", delay_value => 1)  port map(req => inputPort_1_Daemon_CP_3_elements(29), ack => inputPort_1_Daemon_CP_3_elements(31), clk => clk, reset =>reset);
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	57 
    -- CP-element group 32: 	60 
    -- CP-element group 32: 	63 
    -- CP-element group 32: 	66 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_73_update_start_
      -- 
    inputPort_1_Daemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(9) & inputPort_1_Daemon_CP_3_elements(57) & inputPort_1_Daemon_CP_3_elements(60) & inputPort_1_Daemon_CP_3_elements(63) & inputPort_1_Daemon_CP_3_elements(66);
      gj_inputPort_1_Daemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/RPIPE_in_data_1_75_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/RPIPE_in_data_1_75_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/RPIPE_in_data_1_75_Sample/rr
      -- 
    rr_88_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_88_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(33), ack => RPIPE_in_data_1_75_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(11) & inputPort_1_Daemon_CP_3_elements(36);
      gj_inputPort_1_Daemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	13 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/RPIPE_in_data_1_75_update_start_
      -- CP-element group 34: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/RPIPE_in_data_1_75_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/RPIPE_in_data_1_75_Update/cr
      -- 
    cr_93_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_93_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(34), ack => RPIPE_in_data_1_75_inst_req_1); -- 
    inputPort_1_Daemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(13) & inputPort_1_Daemon_CP_3_elements(35);
      gj_inputPort_1_Daemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/RPIPE_in_data_1_75_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/RPIPE_in_data_1_75_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/RPIPE_in_data_1_75_Sample/ra
      -- 
    ra_89_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_1_75_inst_ack_0, ack => inputPort_1_Daemon_CP_3_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	56 
    -- CP-element group 36: 	59 
    -- CP-element group 36: 	62 
    -- CP-element group 36: 	65 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_73_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/RPIPE_in_data_1_75_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/RPIPE_in_data_1_75_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/RPIPE_in_data_1_75_Update/ca
      -- 
    ca_94_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_1_75_inst_ack_1, ack => inputPort_1_Daemon_CP_3_elements(36)); -- 
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	9 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	12 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	11 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_sample_start_
      -- 
    inputPort_1_Daemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(9) & inputPort_1_Daemon_CP_3_elements(12);
      gj_inputPort_1_Daemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	9 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	57 
    -- CP-element group 38: 	60 
    -- CP-element group 38: 	63 
    -- CP-element group 38: 	66 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	13 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_update_start_
      -- 
    inputPort_1_Daemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(9) & inputPort_1_Daemon_CP_3_elements(57) & inputPort_1_Daemon_CP_3_elements(60) & inputPort_1_Daemon_CP_3_elements(63) & inputPort_1_Daemon_CP_3_elements(66);
      gj_inputPort_1_Daemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	11 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_sample_start__ps
      -- 
    inputPort_1_Daemon_CP_3_elements(39) <= inputPort_1_Daemon_CP_3_elements(11);
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	12 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_sample_completed__ps
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	13 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_update_start__ps
      -- 
    inputPort_1_Daemon_CP_3_elements(41) <= inputPort_1_Daemon_CP_3_elements(13);
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	14 
    -- CP-element group 42: 	56 
    -- CP-element group 42: 	59 
    -- CP-element group 42: 	62 
    -- CP-element group 42: 	65 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_update_completed__ps
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	7 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_loopback_trigger
      -- 
    inputPort_1_Daemon_CP_3_elements(43) <= inputPort_1_Daemon_CP_3_elements(7);
    -- CP-element group 44:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_loopback_sample_req
      -- CP-element group 44: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_loopback_sample_req_ps
      -- 
    phi_stmt_76_loopback_sample_req_104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_76_loopback_sample_req_104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(44), ack => phi_stmt_76_req_1); -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	8 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_entry_trigger
      -- 
    inputPort_1_Daemon_CP_3_elements(45) <= inputPort_1_Daemon_CP_3_elements(8);
    -- CP-element group 46:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_entry_sample_req
      -- CP-element group 46: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_entry_sample_req_ps
      -- 
    phi_stmt_76_entry_sample_req_107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_76_entry_sample_req_107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(46), ack => phi_stmt_76_req_0); -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_phi_mux_ack
      -- CP-element group 47: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/phi_stmt_76_phi_mux_ack_ps
      -- 
    phi_stmt_76_phi_mux_ack_110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_76_ack_0, ack => inputPort_1_Daemon_CP_3_elements(47)); -- 
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/konst_78_sample_start__ps
      -- CP-element group 48: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/konst_78_sample_completed__ps
      -- CP-element group 48: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/konst_78_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/konst_78_sample_completed_
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/konst_78_update_start__ps
      -- CP-element group 49: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/konst_78_update_start_
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/konst_78_update_completed__ps
      -- 
    inputPort_1_Daemon_CP_3_elements(50) <= inputPort_1_Daemon_CP_3_elements(51);
    -- CP-element group 51:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	50 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/konst_78_update_completed_
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(51) is a control-delay.
    cp_element_51_delay: control_delay_element  generic map(name => " 51_delay", delay_value => 1)  port map(req => inputPort_1_Daemon_CP_3_elements(49), ack => inputPort_1_Daemon_CP_3_elements(51), clk => clk, reset =>reset);
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_Sample/req
      -- 
    req_131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(52), ack => next_last_dest_id_109_79_buf_req_0); -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_update_start_
      -- CP-element group 53: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_Update/req
      -- 
    req_136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(53), ack => next_last_dest_id_109_79_buf_req_1); -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_Sample/ack
      -- 
    ack_132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_109_79_buf_ack_0, ack => inputPort_1_Daemon_CP_3_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/R_next_last_dest_id_79_Update/ack
      -- 
    ack_137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_109_79_buf_ack_1, ack => inputPort_1_Daemon_CP_3_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	18 
    -- CP-element group 56: 	36 
    -- CP-element group 56: 	42 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_1_121_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_1_121_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_1_121_Sample/req
      -- 
    req_146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(56), ack => WPIPE_noblock_obuf_1_1_121_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(18) & inputPort_1_Daemon_CP_3_elements(36) & inputPort_1_Daemon_CP_3_elements(42) & inputPort_1_Daemon_CP_3_elements(58);
      gj_inputPort_1_Daemon_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	16 
    -- CP-element group 57: 	32 
    -- CP-element group 57: 	38 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_1_121_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_1_121_update_start_
      -- CP-element group 57: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_1_121_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_1_121_Sample/ack
      -- CP-element group 57: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_1_121_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_1_121_Update/req
      -- 
    ack_147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_1_121_inst_ack_0, ack => inputPort_1_Daemon_CP_3_elements(57)); -- 
    req_151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(57), ack => WPIPE_noblock_obuf_1_1_121_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	69 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_1_121_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_1_121_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_1_121_Update/ack
      -- 
    ack_152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_1_121_inst_ack_1, ack => inputPort_1_Daemon_CP_3_elements(58)); -- 
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	18 
    -- CP-element group 59: 	36 
    -- CP-element group 59: 	42 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_2_130_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_2_130_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_2_130_Sample/req
      -- 
    req_160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(59), ack => WPIPE_noblock_obuf_1_2_130_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(18) & inputPort_1_Daemon_CP_3_elements(36) & inputPort_1_Daemon_CP_3_elements(42) & inputPort_1_Daemon_CP_3_elements(61);
      gj_inputPort_1_Daemon_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	16 
    -- CP-element group 60: 	32 
    -- CP-element group 60: 	38 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_2_130_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_2_130_update_start_
      -- CP-element group 60: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_2_130_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_2_130_Sample/ack
      -- CP-element group 60: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_2_130_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_2_130_Update/req
      -- 
    ack_161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_2_130_inst_ack_0, ack => inputPort_1_Daemon_CP_3_elements(60)); -- 
    req_165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(60), ack => WPIPE_noblock_obuf_1_2_130_inst_req_1); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	69 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_2_130_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_2_130_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_2_130_Update/ack
      -- 
    ack_166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_2_130_inst_ack_1, ack => inputPort_1_Daemon_CP_3_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	18 
    -- CP-element group 62: 	36 
    -- CP-element group 62: 	42 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_3_139_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_3_139_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_3_139_Sample/req
      -- 
    req_174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(62), ack => WPIPE_noblock_obuf_1_3_139_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(18) & inputPort_1_Daemon_CP_3_elements(36) & inputPort_1_Daemon_CP_3_elements(42) & inputPort_1_Daemon_CP_3_elements(64);
      gj_inputPort_1_Daemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	16 
    -- CP-element group 63: 	32 
    -- CP-element group 63: 	38 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_3_139_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_3_139_update_start_
      -- CP-element group 63: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_3_139_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_3_139_Sample/ack
      -- CP-element group 63: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_3_139_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_3_139_Update/req
      -- 
    ack_175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_3_139_inst_ack_0, ack => inputPort_1_Daemon_CP_3_elements(63)); -- 
    req_179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(63), ack => WPIPE_noblock_obuf_1_3_139_inst_req_1); -- 
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	69 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_3_139_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_3_139_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_3_139_Update/ack
      -- 
    ack_180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_3_139_inst_ack_1, ack => inputPort_1_Daemon_CP_3_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	18 
    -- CP-element group 65: 	36 
    -- CP-element group 65: 	42 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_4_148_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_4_148_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_4_148_Sample/req
      -- 
    req_188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(65), ack => WPIPE_noblock_obuf_1_4_148_inst_req_0); -- 
    inputPort_1_Daemon_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(18) & inputPort_1_Daemon_CP_3_elements(36) & inputPort_1_Daemon_CP_3_elements(42) & inputPort_1_Daemon_CP_3_elements(67);
      gj_inputPort_1_Daemon_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	16 
    -- CP-element group 66: 	32 
    -- CP-element group 66: 	38 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_4_148_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_4_148_update_start_
      -- CP-element group 66: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_4_148_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_4_148_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_4_148_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_4_148_Update/req
      -- 
    ack_189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_4_148_inst_ack_0, ack => inputPort_1_Daemon_CP_3_elements(66)); -- 
    req_193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_1_Daemon_CP_3_elements(66), ack => WPIPE_noblock_obuf_1_4_148_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_4_148_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_4_148_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/WPIPE_noblock_obuf_1_4_148_Update/ack
      -- 
    ack_194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_1_4_148_inst_ack_1, ack => inputPort_1_Daemon_CP_3_elements(67)); -- 
    -- CP-element group 68:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	9 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	10 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group inputPort_1_Daemon_CP_3_elements(68) is a control-delay.
    cp_element_68_delay: control_delay_element  generic map(name => " 68_delay", delay_value => 1)  port map(req => inputPort_1_Daemon_CP_3_elements(9), ack => inputPort_1_Daemon_CP_3_elements(68), clk => clk, reset =>reset);
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	12 
    -- CP-element group 69: 	58 
    -- CP-element group 69: 	61 
    -- CP-element group 69: 	64 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	6 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_64/do_while_stmt_65/do_while_stmt_65_loop_body/$exit
      -- 
    inputPort_1_Daemon_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_1_Daemon_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_1_Daemon_CP_3_elements(12) & inputPort_1_Daemon_CP_3_elements(58) & inputPort_1_Daemon_CP_3_elements(61) & inputPort_1_Daemon_CP_3_elements(64) & inputPort_1_Daemon_CP_3_elements(67);
      gj_inputPort_1_Daemon_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	5 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_64/do_while_stmt_65/loop_exit/$exit
      -- CP-element group 70: 	 branch_block_stmt_64/do_while_stmt_65/loop_exit/ack
      -- 
    ack_199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_65_branch_ack_0, ack => inputPort_1_Daemon_CP_3_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	5 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_64/do_while_stmt_65/loop_taken/$exit
      -- CP-element group 71: 	 branch_block_stmt_64/do_while_stmt_65/loop_taken/ack
      -- 
    ack_203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_65_branch_ack_1, ack => inputPort_1_Daemon_CP_3_elements(71)); -- 
    -- CP-element group 72:  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	3 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	1 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_64/do_while_stmt_65/$exit
      -- 
    inputPort_1_Daemon_CP_3_elements(72) <= inputPort_1_Daemon_CP_3_elements(3);
    inputPort_1_Daemon_do_while_stmt_65_terminator_204: loop_terminator -- 
      generic map (name => " inputPort_1_Daemon_do_while_stmt_65_terminator_204", max_iterations_in_flight =>7) 
      port map(loop_body_exit => inputPort_1_Daemon_CP_3_elements(6),loop_continue => inputPort_1_Daemon_CP_3_elements(71),loop_terminate => inputPort_1_Daemon_CP_3_elements(70),loop_back => inputPort_1_Daemon_CP_3_elements(4),loop_exit => inputPort_1_Daemon_CP_3_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_67_phi_seq_76_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_1_Daemon_CP_3_elements(19);
      inputPort_1_Daemon_CP_3_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_1_Daemon_CP_3_elements(26);
      inputPort_1_Daemon_CP_3_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_1_Daemon_CP_3_elements(27);
      inputPort_1_Daemon_CP_3_elements(20) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_1_Daemon_CP_3_elements(21);
      inputPort_1_Daemon_CP_3_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_1_Daemon_CP_3_elements(28);
      inputPort_1_Daemon_CP_3_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_1_Daemon_CP_3_elements(30);
      inputPort_1_Daemon_CP_3_elements(22) <= phi_mux_reqs(1);
      phi_stmt_67_phi_seq_76 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_67_phi_seq_76") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_1_Daemon_CP_3_elements(11), 
          phi_sample_ack => inputPort_1_Daemon_CP_3_elements(17), 
          phi_update_req => inputPort_1_Daemon_CP_3_elements(13), 
          phi_update_ack => inputPort_1_Daemon_CP_3_elements(18), 
          phi_mux_ack => inputPort_1_Daemon_CP_3_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_76_phi_seq_138_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_1_Daemon_CP_3_elements(45);
      inputPort_1_Daemon_CP_3_elements(48)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_1_Daemon_CP_3_elements(48);
      inputPort_1_Daemon_CP_3_elements(49)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_1_Daemon_CP_3_elements(50);
      inputPort_1_Daemon_CP_3_elements(46) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_1_Daemon_CP_3_elements(43);
      inputPort_1_Daemon_CP_3_elements(52)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_1_Daemon_CP_3_elements(54);
      inputPort_1_Daemon_CP_3_elements(53)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_1_Daemon_CP_3_elements(55);
      inputPort_1_Daemon_CP_3_elements(44) <= phi_mux_reqs(1);
      phi_stmt_76_phi_seq_138 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_76_phi_seq_138") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_1_Daemon_CP_3_elements(39), 
          phi_sample_ack => inputPort_1_Daemon_CP_3_elements(40), 
          phi_update_req => inputPort_1_Daemon_CP_3_elements(41), 
          phi_update_ack => inputPort_1_Daemon_CP_3_elements(42), 
          phi_mux_ack => inputPort_1_Daemon_CP_3_elements(47), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_28_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= inputPort_1_Daemon_CP_3_elements(7);
        preds(1)  <= inputPort_1_Daemon_CP_3_elements(8);
        entry_tmerge_28 : transition_merge -- 
          generic map(name => " entry_tmerge_28")
          port map (preds => preds, symbol_out => inputPort_1_Daemon_CP_3_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal RPIPE_in_data_1_75_wire : std_logic_vector(31 downto 0);
    signal R_ONE_1_111_wire_constant : std_logic_vector(0 downto 0);
    signal SUB_u16_u16_101_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_98_wire : std_logic_vector(15 downto 0);
    signal count_down_67 : std_logic_vector(15 downto 0);
    signal data_to_outport_114 : std_logic_vector(32 downto 0);
    signal dest_id_89 : std_logic_vector(7 downto 0);
    signal input_word_73 : std_logic_vector(31 downto 0);
    signal konst_100_wire_constant : std_logic_vector(15 downto 0);
    signal konst_117_wire_constant : std_logic_vector(7 downto 0);
    signal konst_126_wire_constant : std_logic_vector(7 downto 0);
    signal konst_135_wire_constant : std_logic_vector(7 downto 0);
    signal konst_144_wire_constant : std_logic_vector(7 downto 0);
    signal konst_152_wire_constant : std_logic_vector(0 downto 0);
    signal konst_78_wire_constant : std_logic_vector(7 downto 0);
    signal konst_83_wire_constant : std_logic_vector(15 downto 0);
    signal konst_97_wire_constant : std_logic_vector(15 downto 0);
    signal last_dest_id_76 : std_logic_vector(7 downto 0);
    signal new_packet_85 : std_logic_vector(0 downto 0);
    signal next_count_down_103 : std_logic_vector(15 downto 0);
    signal next_count_down_103_69_buffered : std_logic_vector(15 downto 0);
    signal next_last_dest_id_109 : std_logic_vector(7 downto 0);
    signal next_last_dest_id_109_79_buffered : std_logic_vector(7 downto 0);
    signal pkt_length_93 : std_logic_vector(15 downto 0);
    signal send_to_1_119 : std_logic_vector(0 downto 0);
    signal send_to_2_128 : std_logic_vector(0 downto 0);
    signal send_to_3_137 : std_logic_vector(0 downto 0);
    signal send_to_4_146 : std_logic_vector(0 downto 0);
    signal type_cast_72_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    R_ONE_1_111_wire_constant <= "1";
    konst_100_wire_constant <= "0000000000000001";
    konst_117_wire_constant <= "00000001";
    konst_126_wire_constant <= "00000010";
    konst_135_wire_constant <= "00000011";
    konst_144_wire_constant <= "00000100";
    konst_152_wire_constant <= "1";
    konst_78_wire_constant <= "00000000";
    konst_83_wire_constant <= "0000000000000000";
    konst_97_wire_constant <= "0000000000000001";
    type_cast_72_wire_constant <= "0000000000000000";
    phi_stmt_67: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= next_count_down_103_69_buffered & type_cast_72_wire_constant;
      req <= phi_stmt_67_req_0 & phi_stmt_67_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_67",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_67_ack_0,
          idata => idata,
          odata => count_down_67,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_67
    phi_stmt_76: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_78_wire_constant & next_last_dest_id_109_79_buffered;
      req <= phi_stmt_76_req_0 & phi_stmt_76_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_76",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_76_ack_0,
          idata => idata,
          odata => last_dest_id_76,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_76
    -- flow-through select operator MUX_102_inst
    next_count_down_103 <= SUB_u16_u16_98_wire when (new_packet_85(0) /=  '0') else SUB_u16_u16_101_wire;
    -- flow-through select operator MUX_108_inst
    next_last_dest_id_109 <= dest_id_89 when (new_packet_85(0) /=  '0') else last_dest_id_76;
    -- flow-through slice operator slice_88_inst
    dest_id_89 <= input_word_73(31 downto 24);
    -- flow-through slice operator slice_92_inst
    pkt_length_93 <= input_word_73(23 downto 8);
    next_count_down_103_69_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_count_down_103_69_buf_req_0;
      next_count_down_103_69_buf_ack_0<= wack(0);
      rreq(0) <= next_count_down_103_69_buf_req_1;
      next_count_down_103_69_buf_ack_1<= rack(0);
      next_count_down_103_69_buf : InterlockBuffer generic map ( -- 
        name => "next_count_down_103_69_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_count_down_103,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_count_down_103_69_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_last_dest_id_109_79_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_last_dest_id_109_79_buf_req_0;
      next_last_dest_id_109_79_buf_ack_0<= wack(0);
      rreq(0) <= next_last_dest_id_109_79_buf_req_1;
      next_last_dest_id_109_79_buf_ack_1<= rack(0);
      next_last_dest_id_109_79_buf : InterlockBuffer generic map ( -- 
        name => "next_last_dest_id_109_79_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_last_dest_id_109,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_last_dest_id_109_79_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_73
    process(RPIPE_in_data_1_75_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := RPIPE_in_data_1_75_wire(31 downto 0);
      input_word_73 <= tmp_var; -- 
    end process;
    do_while_stmt_65_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_152_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_65_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_65_branch_req_0,
          ack0 => do_while_stmt_65_branch_ack_0,
          ack1 => do_while_stmt_65_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator CONCAT_u1_u33_113_inst
    process(R_ONE_1_111_wire_constant, input_word_73) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ONE_1_111_wire_constant, input_word_73, tmp_var);
      data_to_outport_114 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_84_inst
    process(count_down_67) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(count_down_67, konst_83_wire_constant, tmp_var);
      new_packet_85 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_118_inst
    process(next_last_dest_id_109) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_109, konst_117_wire_constant, tmp_var);
      send_to_1_119 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_127_inst
    process(next_last_dest_id_109) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_109, konst_126_wire_constant, tmp_var);
      send_to_2_128 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_136_inst
    process(next_last_dest_id_109) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_109, konst_135_wire_constant, tmp_var);
      send_to_3_137 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_145_inst
    process(next_last_dest_id_109) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_109, konst_144_wire_constant, tmp_var);
      send_to_4_146 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_101_inst
    process(count_down_67) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(count_down_67, konst_100_wire_constant, tmp_var);
      SUB_u16_u16_101_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_98_inst
    process(pkt_length_93) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(pkt_length_93, konst_97_wire_constant, tmp_var);
      SUB_u16_u16_98_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_in_data_1_75_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_in_data_1_75_inst_req_0;
      RPIPE_in_data_1_75_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_in_data_1_75_inst_req_1;
      RPIPE_in_data_1_75_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_in_data_1_75_wire <= data_out(31 downto 0);
      in_data_1_read_0_gI: SplitGuardInterface generic map(name => "in_data_1_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      in_data_1_read_0: InputPortRevised -- 
        generic map ( name => "in_data_1_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => in_data_1_pipe_read_req(0),
          oack => in_data_1_pipe_read_ack(0),
          odata => in_data_1_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_noblock_obuf_1_1_121_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_1_1_121_inst_req_0;
      WPIPE_noblock_obuf_1_1_121_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_1_1_121_inst_req_1;
      WPIPE_noblock_obuf_1_1_121_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_1_119(0);
      data_in <= data_to_outport_114;
      noblock_obuf_1_1_write_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_1_write_0: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_1_1", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_1_1_pipe_write_req(0),
          oack => noblock_obuf_1_1_pipe_write_ack(0),
          odata => noblock_obuf_1_1_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_noblock_obuf_1_2_130_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_1_2_130_inst_req_0;
      WPIPE_noblock_obuf_1_2_130_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_1_2_130_inst_req_1;
      WPIPE_noblock_obuf_1_2_130_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_2_128(0);
      data_in <= data_to_outport_114;
      noblock_obuf_1_2_write_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_2_write_1: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_1_2", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_1_2_pipe_write_req(0),
          oack => noblock_obuf_1_2_pipe_write_ack(0),
          odata => noblock_obuf_1_2_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_noblock_obuf_1_3_139_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_1_3_139_inst_req_0;
      WPIPE_noblock_obuf_1_3_139_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_1_3_139_inst_req_1;
      WPIPE_noblock_obuf_1_3_139_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_3_137(0);
      data_in <= data_to_outport_114;
      noblock_obuf_1_3_write_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_3_write_2: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_1_3", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_1_3_pipe_write_req(0),
          oack => noblock_obuf_1_3_pipe_write_ack(0),
          odata => noblock_obuf_1_3_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_noblock_obuf_1_4_148_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_1_4_148_inst_req_0;
      WPIPE_noblock_obuf_1_4_148_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_1_4_148_inst_req_1;
      WPIPE_noblock_obuf_1_4_148_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_4_146(0);
      data_in <= data_to_outport_114;
      noblock_obuf_1_4_write_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_4_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_4_write_3: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_1_4", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_1_4_pipe_write_req(0),
          oack => noblock_obuf_1_4_pipe_write_ack(0),
          odata => noblock_obuf_1_4_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end inputPort_1_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity inputPort_2_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    in_data_2_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_2_pipe_read_data : in   std_logic_vector(31 downto 0);
    noblock_obuf_2_1_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_1_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_2_2_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_2_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_2_3_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_3_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_2_4_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_4_pipe_write_data : out  std_logic_vector(32 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity inputPort_2_Daemon;
architecture inputPort_2_Daemon_arch of inputPort_2_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal inputPort_2_Daemon_CP_205_start: Boolean;
  signal inputPort_2_Daemon_CP_205_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_noblock_obuf_2_3_230_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_2_3_230_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_2_3_230_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_2_3_230_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_2_4_239_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_2_4_239_inst_ack_0 : boolean;
  signal do_while_stmt_157_branch_req_0 : boolean;
  signal phi_stmt_159_req_0 : boolean;
  signal phi_stmt_159_req_1 : boolean;
  signal phi_stmt_159_ack_0 : boolean;
  signal next_count_down_194_161_buf_req_0 : boolean;
  signal next_count_down_194_161_buf_ack_0 : boolean;
  signal next_count_down_194_161_buf_req_1 : boolean;
  signal next_count_down_194_161_buf_ack_1 : boolean;
  signal RPIPE_in_data_2_166_inst_req_0 : boolean;
  signal RPIPE_in_data_2_166_inst_ack_0 : boolean;
  signal RPIPE_in_data_2_166_inst_req_1 : boolean;
  signal RPIPE_in_data_2_166_inst_ack_1 : boolean;
  signal phi_stmt_167_req_1 : boolean;
  signal phi_stmt_167_req_0 : boolean;
  signal phi_stmt_167_ack_0 : boolean;
  signal next_last_dest_id_200_170_buf_req_0 : boolean;
  signal next_last_dest_id_200_170_buf_ack_0 : boolean;
  signal next_last_dest_id_200_170_buf_req_1 : boolean;
  signal next_last_dest_id_200_170_buf_ack_1 : boolean;
  signal WPIPE_noblock_obuf_2_1_212_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_2_1_212_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_2_1_212_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_2_1_212_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_2_2_221_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_2_2_221_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_2_2_221_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_2_2_221_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_2_4_239_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_2_4_239_inst_ack_1 : boolean;
  signal do_while_stmt_157_branch_ack_0 : boolean;
  signal do_while_stmt_157_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "inputPort_2_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  inputPort_2_Daemon_CP_205_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "inputPort_2_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_2_Daemon_CP_205_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= inputPort_2_Daemon_CP_205_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_2_Daemon_CP_205_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  inputPort_2_Daemon_CP_205: Block -- control-path 
    signal inputPort_2_Daemon_CP_205_elements: BooleanArray(72 downto 0);
    -- 
  begin -- 
    inputPort_2_Daemon_CP_205_elements(0) <= inputPort_2_Daemon_CP_205_start;
    inputPort_2_Daemon_CP_205_symbol <= inputPort_2_Daemon_CP_205_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_156/$entry
      -- CP-element group 0: 	 branch_block_stmt_156/branch_block_stmt_156__entry__
      -- CP-element group 0: 	 branch_block_stmt_156/do_while_stmt_157__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	72 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_156/$exit
      -- CP-element group 1: 	 branch_block_stmt_156/branch_block_stmt_156__exit__
      -- CP-element group 1: 	 branch_block_stmt_156/do_while_stmt_157__exit__
      -- 
    inputPort_2_Daemon_CP_205_elements(1) <= inputPort_2_Daemon_CP_205_elements(72);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_156/do_while_stmt_157/$entry
      -- CP-element group 2: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157__entry__
      -- 
    inputPort_2_Daemon_CP_205_elements(2) <= inputPort_2_Daemon_CP_205_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	72 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157__exit__
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_156/do_while_stmt_157/loop_back
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	70 
    -- CP-element group 5: 	71 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_156/do_while_stmt_157/condition_done
      -- CP-element group 5: 	 branch_block_stmt_156/do_while_stmt_157/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_156/do_while_stmt_157/loop_taken/$entry
      -- 
    inputPort_2_Daemon_CP_205_elements(5) <= inputPort_2_Daemon_CP_205_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	69 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_156/do_while_stmt_157/loop_body_done
      -- 
    inputPort_2_Daemon_CP_205_elements(6) <= inputPort_2_Daemon_CP_205_elements(69);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	43 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/back_edge_to_loop_body
      -- 
    inputPort_2_Daemon_CP_205_elements(7) <= inputPort_2_Daemon_CP_205_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	45 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/first_time_through_loop_body
      -- 
    inputPort_2_Daemon_CP_205_elements(8) <= inputPort_2_Daemon_CP_205_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	37 
    -- CP-element group 9: 	38 
    -- CP-element group 9: 	68 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_164_sample_start_
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	68 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/condition_evaluated
      -- 
    condition_evaluated_229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(10), ack => do_while_stmt_157_branch_req_0); -- 
    inputPort_2_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(14) & inputPort_2_Daemon_CP_205_elements(68);
      gj_inputPort_2_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	37 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11: 	39 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_sample_start__ps
      -- 
    inputPort_2_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(9) & inputPort_2_Daemon_CP_205_elements(15) & inputPort_2_Daemon_CP_205_elements(37) & inputPort_2_Daemon_CP_205_elements(14);
      gj_inputPort_2_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	40 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	69 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	37 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_164_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_sample_completed_
      -- 
    inputPort_2_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(17) & inputPort_2_Daemon_CP_205_elements(35) & inputPort_2_Daemon_CP_205_elements(40);
      gj_inputPort_2_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	32 
    -- CP-element group 13: 	38 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13: 	41 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_update_start__ps
      -- 
    inputPort_2_Daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(16) & inputPort_2_Daemon_CP_205_elements(32) & inputPort_2_Daemon_CP_205_elements(38);
      gj_inputPort_2_Daemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	36 
    -- CP-element group 14: 	42 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/aggregated_phi_update_ack
      -- 
    inputPort_2_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(18) & inputPort_2_Daemon_CP_205_elements(36) & inputPort_2_Daemon_CP_205_elements(42);
      gj_inputPort_2_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_sample_start_
      -- 
    inputPort_2_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(9) & inputPort_2_Daemon_CP_205_elements(12);
      gj_inputPort_2_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	57 
    -- CP-element group 16: 	60 
    -- CP-element group 16: 	63 
    -- CP-element group 16: 	66 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_update_start_
      -- 
    inputPort_2_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(9) & inputPort_2_Daemon_CP_205_elements(57) & inputPort_2_Daemon_CP_205_elements(60) & inputPort_2_Daemon_CP_205_elements(63) & inputPort_2_Daemon_CP_205_elements(66);
      gj_inputPort_2_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_sample_completed__ps
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	56 
    -- CP-element group 18: 	59 
    -- CP-element group 18: 	62 
    -- CP-element group 18: 	65 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_update_completed__ps
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_loopback_trigger
      -- 
    inputPort_2_Daemon_CP_205_elements(19) <= inputPort_2_Daemon_CP_205_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_loopback_sample_req_ps
      -- 
    phi_stmt_159_loopback_sample_req_244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_159_loopback_sample_req_244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(20), ack => phi_stmt_159_req_0); -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_entry_trigger
      -- 
    inputPort_2_Daemon_CP_205_elements(21) <= inputPort_2_Daemon_CP_205_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_entry_sample_req_ps
      -- 
    phi_stmt_159_entry_sample_req_247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_159_entry_sample_req_247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(22), ack => phi_stmt_159_req_1); -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_159_phi_mux_ack_ps
      -- 
    phi_stmt_159_phi_mux_ack_250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_159_ack_0, ack => inputPort_2_Daemon_CP_205_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_Sample/req
      -- 
    req_263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(24), ack => next_count_down_194_161_buf_req_0); -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_update_start_
      -- CP-element group 25: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_Update/req
      -- 
    req_268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(25), ack => next_count_down_194_161_buf_req_1); -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_Sample/ack
      -- 
    ack_264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_194_161_buf_ack_0, ack => inputPort_2_Daemon_CP_205_elements(26)); -- 
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_update_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_count_down_161_Update/ack
      -- 
    ack_269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_194_161_buf_ack_1, ack => inputPort_2_Daemon_CP_205_elements(27)); -- 
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/type_cast_163_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/type_cast_163_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/type_cast_163_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/type_cast_163_sample_completed_
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/type_cast_163_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/type_cast_163_update_start_
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/type_cast_163_update_completed__ps
      -- 
    inputPort_2_Daemon_CP_205_elements(30) <= inputPort_2_Daemon_CP_205_elements(31);
    -- CP-element group 31:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	30 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/type_cast_163_update_completed_
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(31) is a control-delay.
    cp_element_31_delay: control_delay_element  generic map(name => " 31_delay", delay_value => 1)  port map(req => inputPort_2_Daemon_CP_205_elements(29), ack => inputPort_2_Daemon_CP_205_elements(31), clk => clk, reset =>reset);
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	57 
    -- CP-element group 32: 	60 
    -- CP-element group 32: 	63 
    -- CP-element group 32: 	66 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_164_update_start_
      -- 
    inputPort_2_Daemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(9) & inputPort_2_Daemon_CP_205_elements(57) & inputPort_2_Daemon_CP_205_elements(60) & inputPort_2_Daemon_CP_205_elements(63) & inputPort_2_Daemon_CP_205_elements(66);
      gj_inputPort_2_Daemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/RPIPE_in_data_2_166_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/RPIPE_in_data_2_166_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/RPIPE_in_data_2_166_Sample/rr
      -- 
    rr_290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(33), ack => RPIPE_in_data_2_166_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(11) & inputPort_2_Daemon_CP_205_elements(36);
      gj_inputPort_2_Daemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	13 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/RPIPE_in_data_2_166_update_start_
      -- CP-element group 34: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/RPIPE_in_data_2_166_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/RPIPE_in_data_2_166_Update/cr
      -- 
    cr_295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(34), ack => RPIPE_in_data_2_166_inst_req_1); -- 
    inputPort_2_Daemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(13) & inputPort_2_Daemon_CP_205_elements(35);
      gj_inputPort_2_Daemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/RPIPE_in_data_2_166_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/RPIPE_in_data_2_166_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/RPIPE_in_data_2_166_Sample/ra
      -- 
    ra_291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_2_166_inst_ack_0, ack => inputPort_2_Daemon_CP_205_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	56 
    -- CP-element group 36: 	59 
    -- CP-element group 36: 	62 
    -- CP-element group 36: 	65 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_164_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/RPIPE_in_data_2_166_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/RPIPE_in_data_2_166_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/RPIPE_in_data_2_166_Update/ca
      -- 
    ca_296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_2_166_inst_ack_1, ack => inputPort_2_Daemon_CP_205_elements(36)); -- 
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	9 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	12 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	11 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_sample_start_
      -- 
    inputPort_2_Daemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(9) & inputPort_2_Daemon_CP_205_elements(12);
      gj_inputPort_2_Daemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	9 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	57 
    -- CP-element group 38: 	60 
    -- CP-element group 38: 	63 
    -- CP-element group 38: 	66 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	13 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_update_start_
      -- 
    inputPort_2_Daemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(9) & inputPort_2_Daemon_CP_205_elements(57) & inputPort_2_Daemon_CP_205_elements(60) & inputPort_2_Daemon_CP_205_elements(63) & inputPort_2_Daemon_CP_205_elements(66);
      gj_inputPort_2_Daemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	11 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_sample_start__ps
      -- 
    inputPort_2_Daemon_CP_205_elements(39) <= inputPort_2_Daemon_CP_205_elements(11);
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	12 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_sample_completed__ps
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	13 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_update_start__ps
      -- 
    inputPort_2_Daemon_CP_205_elements(41) <= inputPort_2_Daemon_CP_205_elements(13);
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	14 
    -- CP-element group 42: 	56 
    -- CP-element group 42: 	59 
    -- CP-element group 42: 	62 
    -- CP-element group 42: 	65 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_update_completed__ps
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	7 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_loopback_trigger
      -- 
    inputPort_2_Daemon_CP_205_elements(43) <= inputPort_2_Daemon_CP_205_elements(7);
    -- CP-element group 44:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_loopback_sample_req
      -- CP-element group 44: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_loopback_sample_req_ps
      -- 
    phi_stmt_167_loopback_sample_req_306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_167_loopback_sample_req_306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(44), ack => phi_stmt_167_req_1); -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	8 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_entry_trigger
      -- 
    inputPort_2_Daemon_CP_205_elements(45) <= inputPort_2_Daemon_CP_205_elements(8);
    -- CP-element group 46:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_entry_sample_req
      -- CP-element group 46: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_entry_sample_req_ps
      -- 
    phi_stmt_167_entry_sample_req_309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_167_entry_sample_req_309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(46), ack => phi_stmt_167_req_0); -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_phi_mux_ack
      -- CP-element group 47: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/phi_stmt_167_phi_mux_ack_ps
      -- 
    phi_stmt_167_phi_mux_ack_312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_167_ack_0, ack => inputPort_2_Daemon_CP_205_elements(47)); -- 
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/konst_169_sample_start__ps
      -- CP-element group 48: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/konst_169_sample_completed__ps
      -- CP-element group 48: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/konst_169_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/konst_169_sample_completed_
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/konst_169_update_start__ps
      -- CP-element group 49: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/konst_169_update_start_
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/konst_169_update_completed__ps
      -- 
    inputPort_2_Daemon_CP_205_elements(50) <= inputPort_2_Daemon_CP_205_elements(51);
    -- CP-element group 51:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	50 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/konst_169_update_completed_
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(51) is a control-delay.
    cp_element_51_delay: control_delay_element  generic map(name => " 51_delay", delay_value => 1)  port map(req => inputPort_2_Daemon_CP_205_elements(49), ack => inputPort_2_Daemon_CP_205_elements(51), clk => clk, reset =>reset);
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_Sample/req
      -- 
    req_333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(52), ack => next_last_dest_id_200_170_buf_req_0); -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_update_start_
      -- CP-element group 53: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_Update/req
      -- 
    req_338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(53), ack => next_last_dest_id_200_170_buf_req_1); -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_Sample/ack
      -- 
    ack_334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_200_170_buf_ack_0, ack => inputPort_2_Daemon_CP_205_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/R_next_last_dest_id_170_Update/ack
      -- 
    ack_339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_200_170_buf_ack_1, ack => inputPort_2_Daemon_CP_205_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	18 
    -- CP-element group 56: 	36 
    -- CP-element group 56: 	42 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_1_212_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_1_212_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_1_212_Sample/req
      -- 
    req_348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(56), ack => WPIPE_noblock_obuf_2_1_212_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(18) & inputPort_2_Daemon_CP_205_elements(36) & inputPort_2_Daemon_CP_205_elements(42) & inputPort_2_Daemon_CP_205_elements(58);
      gj_inputPort_2_Daemon_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	16 
    -- CP-element group 57: 	32 
    -- CP-element group 57: 	38 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_1_212_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_1_212_update_start_
      -- CP-element group 57: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_1_212_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_1_212_Sample/ack
      -- CP-element group 57: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_1_212_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_1_212_Update/req
      -- 
    ack_349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_1_212_inst_ack_0, ack => inputPort_2_Daemon_CP_205_elements(57)); -- 
    req_353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(57), ack => WPIPE_noblock_obuf_2_1_212_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	69 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_1_212_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_1_212_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_1_212_Update/ack
      -- 
    ack_354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_1_212_inst_ack_1, ack => inputPort_2_Daemon_CP_205_elements(58)); -- 
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	18 
    -- CP-element group 59: 	36 
    -- CP-element group 59: 	42 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_2_221_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_2_221_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_2_221_Sample/req
      -- 
    req_362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(59), ack => WPIPE_noblock_obuf_2_2_221_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(18) & inputPort_2_Daemon_CP_205_elements(36) & inputPort_2_Daemon_CP_205_elements(42) & inputPort_2_Daemon_CP_205_elements(61);
      gj_inputPort_2_Daemon_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	16 
    -- CP-element group 60: 	32 
    -- CP-element group 60: 	38 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_2_221_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_2_221_update_start_
      -- CP-element group 60: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_2_221_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_2_221_Sample/ack
      -- CP-element group 60: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_2_221_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_2_221_Update/req
      -- 
    ack_363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_2_221_inst_ack_0, ack => inputPort_2_Daemon_CP_205_elements(60)); -- 
    req_367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(60), ack => WPIPE_noblock_obuf_2_2_221_inst_req_1); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	69 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_2_221_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_2_221_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_2_221_Update/ack
      -- 
    ack_368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_2_221_inst_ack_1, ack => inputPort_2_Daemon_CP_205_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	18 
    -- CP-element group 62: 	36 
    -- CP-element group 62: 	42 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_3_230_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_3_230_Sample/req
      -- CP-element group 62: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_3_230_sample_start_
      -- 
    req_376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(62), ack => WPIPE_noblock_obuf_2_3_230_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(18) & inputPort_2_Daemon_CP_205_elements(36) & inputPort_2_Daemon_CP_205_elements(42) & inputPort_2_Daemon_CP_205_elements(64);
      gj_inputPort_2_Daemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	16 
    -- CP-element group 63: 	32 
    -- CP-element group 63: 	38 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_3_230_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_3_230_Sample/ack
      -- CP-element group 63: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_3_230_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_3_230_Update/req
      -- CP-element group 63: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_3_230_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_3_230_update_start_
      -- 
    ack_377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_3_230_inst_ack_0, ack => inputPort_2_Daemon_CP_205_elements(63)); -- 
    req_381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(63), ack => WPIPE_noblock_obuf_2_3_230_inst_req_1); -- 
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	69 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_3_230_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_3_230_Update/ack
      -- CP-element group 64: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_3_230_update_completed_
      -- 
    ack_382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_3_230_inst_ack_1, ack => inputPort_2_Daemon_CP_205_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	18 
    -- CP-element group 65: 	36 
    -- CP-element group 65: 	42 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_4_239_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_4_239_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_4_239_Sample/req
      -- 
    req_390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(65), ack => WPIPE_noblock_obuf_2_4_239_inst_req_0); -- 
    inputPort_2_Daemon_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(18) & inputPort_2_Daemon_CP_205_elements(36) & inputPort_2_Daemon_CP_205_elements(42) & inputPort_2_Daemon_CP_205_elements(67);
      gj_inputPort_2_Daemon_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	16 
    -- CP-element group 66: 	32 
    -- CP-element group 66: 	38 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_4_239_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_4_239_update_start_
      -- CP-element group 66: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_4_239_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_4_239_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_4_239_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_4_239_Update/req
      -- 
    ack_391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_4_239_inst_ack_0, ack => inputPort_2_Daemon_CP_205_elements(66)); -- 
    req_395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_2_Daemon_CP_205_elements(66), ack => WPIPE_noblock_obuf_2_4_239_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_4_239_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_4_239_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/WPIPE_noblock_obuf_2_4_239_Update/ack
      -- 
    ack_396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_2_4_239_inst_ack_1, ack => inputPort_2_Daemon_CP_205_elements(67)); -- 
    -- CP-element group 68:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	9 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	10 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group inputPort_2_Daemon_CP_205_elements(68) is a control-delay.
    cp_element_68_delay: control_delay_element  generic map(name => " 68_delay", delay_value => 1)  port map(req => inputPort_2_Daemon_CP_205_elements(9), ack => inputPort_2_Daemon_CP_205_elements(68), clk => clk, reset =>reset);
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	12 
    -- CP-element group 69: 	58 
    -- CP-element group 69: 	61 
    -- CP-element group 69: 	64 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	6 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_156/do_while_stmt_157/do_while_stmt_157_loop_body/$exit
      -- 
    inputPort_2_Daemon_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_2_Daemon_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_2_Daemon_CP_205_elements(12) & inputPort_2_Daemon_CP_205_elements(58) & inputPort_2_Daemon_CP_205_elements(61) & inputPort_2_Daemon_CP_205_elements(64) & inputPort_2_Daemon_CP_205_elements(67);
      gj_inputPort_2_Daemon_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	5 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_156/do_while_stmt_157/loop_exit/$exit
      -- CP-element group 70: 	 branch_block_stmt_156/do_while_stmt_157/loop_exit/ack
      -- 
    ack_401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_157_branch_ack_0, ack => inputPort_2_Daemon_CP_205_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	5 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_156/do_while_stmt_157/loop_taken/$exit
      -- CP-element group 71: 	 branch_block_stmt_156/do_while_stmt_157/loop_taken/ack
      -- 
    ack_405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_157_branch_ack_1, ack => inputPort_2_Daemon_CP_205_elements(71)); -- 
    -- CP-element group 72:  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	3 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	1 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_156/do_while_stmt_157/$exit
      -- 
    inputPort_2_Daemon_CP_205_elements(72) <= inputPort_2_Daemon_CP_205_elements(3);
    inputPort_2_Daemon_do_while_stmt_157_terminator_406: loop_terminator -- 
      generic map (name => " inputPort_2_Daemon_do_while_stmt_157_terminator_406", max_iterations_in_flight =>7) 
      port map(loop_body_exit => inputPort_2_Daemon_CP_205_elements(6),loop_continue => inputPort_2_Daemon_CP_205_elements(71),loop_terminate => inputPort_2_Daemon_CP_205_elements(70),loop_back => inputPort_2_Daemon_CP_205_elements(4),loop_exit => inputPort_2_Daemon_CP_205_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_159_phi_seq_278_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_2_Daemon_CP_205_elements(19);
      inputPort_2_Daemon_CP_205_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_2_Daemon_CP_205_elements(26);
      inputPort_2_Daemon_CP_205_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_2_Daemon_CP_205_elements(27);
      inputPort_2_Daemon_CP_205_elements(20) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_2_Daemon_CP_205_elements(21);
      inputPort_2_Daemon_CP_205_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_2_Daemon_CP_205_elements(28);
      inputPort_2_Daemon_CP_205_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_2_Daemon_CP_205_elements(30);
      inputPort_2_Daemon_CP_205_elements(22) <= phi_mux_reqs(1);
      phi_stmt_159_phi_seq_278 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_159_phi_seq_278") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_2_Daemon_CP_205_elements(11), 
          phi_sample_ack => inputPort_2_Daemon_CP_205_elements(17), 
          phi_update_req => inputPort_2_Daemon_CP_205_elements(13), 
          phi_update_ack => inputPort_2_Daemon_CP_205_elements(18), 
          phi_mux_ack => inputPort_2_Daemon_CP_205_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_167_phi_seq_340_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_2_Daemon_CP_205_elements(45);
      inputPort_2_Daemon_CP_205_elements(48)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_2_Daemon_CP_205_elements(48);
      inputPort_2_Daemon_CP_205_elements(49)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_2_Daemon_CP_205_elements(50);
      inputPort_2_Daemon_CP_205_elements(46) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_2_Daemon_CP_205_elements(43);
      inputPort_2_Daemon_CP_205_elements(52)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_2_Daemon_CP_205_elements(54);
      inputPort_2_Daemon_CP_205_elements(53)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_2_Daemon_CP_205_elements(55);
      inputPort_2_Daemon_CP_205_elements(44) <= phi_mux_reqs(1);
      phi_stmt_167_phi_seq_340 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_167_phi_seq_340") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_2_Daemon_CP_205_elements(39), 
          phi_sample_ack => inputPort_2_Daemon_CP_205_elements(40), 
          phi_update_req => inputPort_2_Daemon_CP_205_elements(41), 
          phi_update_ack => inputPort_2_Daemon_CP_205_elements(42), 
          phi_mux_ack => inputPort_2_Daemon_CP_205_elements(47), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_230_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= inputPort_2_Daemon_CP_205_elements(7);
        preds(1)  <= inputPort_2_Daemon_CP_205_elements(8);
        entry_tmerge_230 : transition_merge -- 
          generic map(name => " entry_tmerge_230")
          port map (preds => preds, symbol_out => inputPort_2_Daemon_CP_205_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal RPIPE_in_data_2_166_wire : std_logic_vector(31 downto 0);
    signal R_ONE_1_202_wire_constant : std_logic_vector(0 downto 0);
    signal SUB_u16_u16_189_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_192_wire : std_logic_vector(15 downto 0);
    signal count_down_159 : std_logic_vector(15 downto 0);
    signal data_to_outport_205 : std_logic_vector(32 downto 0);
    signal dest_id_180 : std_logic_vector(7 downto 0);
    signal input_word_164 : std_logic_vector(31 downto 0);
    signal konst_169_wire_constant : std_logic_vector(7 downto 0);
    signal konst_174_wire_constant : std_logic_vector(15 downto 0);
    signal konst_188_wire_constant : std_logic_vector(15 downto 0);
    signal konst_191_wire_constant : std_logic_vector(15 downto 0);
    signal konst_208_wire_constant : std_logic_vector(7 downto 0);
    signal konst_217_wire_constant : std_logic_vector(7 downto 0);
    signal konst_226_wire_constant : std_logic_vector(7 downto 0);
    signal konst_235_wire_constant : std_logic_vector(7 downto 0);
    signal konst_243_wire_constant : std_logic_vector(0 downto 0);
    signal last_dest_id_167 : std_logic_vector(7 downto 0);
    signal new_packet_176 : std_logic_vector(0 downto 0);
    signal next_count_down_194 : std_logic_vector(15 downto 0);
    signal next_count_down_194_161_buffered : std_logic_vector(15 downto 0);
    signal next_last_dest_id_200 : std_logic_vector(7 downto 0);
    signal next_last_dest_id_200_170_buffered : std_logic_vector(7 downto 0);
    signal pkt_length_184 : std_logic_vector(15 downto 0);
    signal send_to_1_210 : std_logic_vector(0 downto 0);
    signal send_to_2_219 : std_logic_vector(0 downto 0);
    signal send_to_3_228 : std_logic_vector(0 downto 0);
    signal send_to_4_237 : std_logic_vector(0 downto 0);
    signal type_cast_163_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    R_ONE_1_202_wire_constant <= "1";
    konst_169_wire_constant <= "00000000";
    konst_174_wire_constant <= "0000000000000000";
    konst_188_wire_constant <= "0000000000000001";
    konst_191_wire_constant <= "0000000000000001";
    konst_208_wire_constant <= "00000001";
    konst_217_wire_constant <= "00000010";
    konst_226_wire_constant <= "00000011";
    konst_235_wire_constant <= "00000100";
    konst_243_wire_constant <= "1";
    type_cast_163_wire_constant <= "0000000000000000";
    phi_stmt_159: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= next_count_down_194_161_buffered & type_cast_163_wire_constant;
      req <= phi_stmt_159_req_0 & phi_stmt_159_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_159",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_159_ack_0,
          idata => idata,
          odata => count_down_159,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_159
    phi_stmt_167: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_169_wire_constant & next_last_dest_id_200_170_buffered;
      req <= phi_stmt_167_req_0 & phi_stmt_167_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_167",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_167_ack_0,
          idata => idata,
          odata => last_dest_id_167,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_167
    -- flow-through select operator MUX_193_inst
    next_count_down_194 <= SUB_u16_u16_189_wire when (new_packet_176(0) /=  '0') else SUB_u16_u16_192_wire;
    -- flow-through select operator MUX_199_inst
    next_last_dest_id_200 <= dest_id_180 when (new_packet_176(0) /=  '0') else last_dest_id_167;
    -- flow-through slice operator slice_179_inst
    dest_id_180 <= input_word_164(31 downto 24);
    -- flow-through slice operator slice_183_inst
    pkt_length_184 <= input_word_164(23 downto 8);
    next_count_down_194_161_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_count_down_194_161_buf_req_0;
      next_count_down_194_161_buf_ack_0<= wack(0);
      rreq(0) <= next_count_down_194_161_buf_req_1;
      next_count_down_194_161_buf_ack_1<= rack(0);
      next_count_down_194_161_buf : InterlockBuffer generic map ( -- 
        name => "next_count_down_194_161_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_count_down_194,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_count_down_194_161_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_last_dest_id_200_170_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_last_dest_id_200_170_buf_req_0;
      next_last_dest_id_200_170_buf_ack_0<= wack(0);
      rreq(0) <= next_last_dest_id_200_170_buf_req_1;
      next_last_dest_id_200_170_buf_ack_1<= rack(0);
      next_last_dest_id_200_170_buf : InterlockBuffer generic map ( -- 
        name => "next_last_dest_id_200_170_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_last_dest_id_200,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_last_dest_id_200_170_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_164
    process(RPIPE_in_data_2_166_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := RPIPE_in_data_2_166_wire(31 downto 0);
      input_word_164 <= tmp_var; -- 
    end process;
    do_while_stmt_157_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_243_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_157_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_157_branch_req_0,
          ack0 => do_while_stmt_157_branch_ack_0,
          ack1 => do_while_stmt_157_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator CONCAT_u1_u33_204_inst
    process(R_ONE_1_202_wire_constant, input_word_164) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ONE_1_202_wire_constant, input_word_164, tmp_var);
      data_to_outport_205 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_175_inst
    process(count_down_159) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(count_down_159, konst_174_wire_constant, tmp_var);
      new_packet_176 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_209_inst
    process(next_last_dest_id_200) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_200, konst_208_wire_constant, tmp_var);
      send_to_1_210 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_218_inst
    process(next_last_dest_id_200) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_200, konst_217_wire_constant, tmp_var);
      send_to_2_219 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_227_inst
    process(next_last_dest_id_200) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_200, konst_226_wire_constant, tmp_var);
      send_to_3_228 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_236_inst
    process(next_last_dest_id_200) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_200, konst_235_wire_constant, tmp_var);
      send_to_4_237 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_189_inst
    process(pkt_length_184) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(pkt_length_184, konst_188_wire_constant, tmp_var);
      SUB_u16_u16_189_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_192_inst
    process(count_down_159) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(count_down_159, konst_191_wire_constant, tmp_var);
      SUB_u16_u16_192_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_in_data_2_166_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_in_data_2_166_inst_req_0;
      RPIPE_in_data_2_166_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_in_data_2_166_inst_req_1;
      RPIPE_in_data_2_166_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_in_data_2_166_wire <= data_out(31 downto 0);
      in_data_2_read_0_gI: SplitGuardInterface generic map(name => "in_data_2_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      in_data_2_read_0: InputPortRevised -- 
        generic map ( name => "in_data_2_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => in_data_2_pipe_read_req(0),
          oack => in_data_2_pipe_read_ack(0),
          odata => in_data_2_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_noblock_obuf_2_1_212_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_2_1_212_inst_req_0;
      WPIPE_noblock_obuf_2_1_212_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_2_1_212_inst_req_1;
      WPIPE_noblock_obuf_2_1_212_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_1_210(0);
      data_in <= data_to_outport_205;
      noblock_obuf_2_1_write_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_1_write_0: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_2_1", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_2_1_pipe_write_req(0),
          oack => noblock_obuf_2_1_pipe_write_ack(0),
          odata => noblock_obuf_2_1_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_noblock_obuf_2_2_221_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_2_2_221_inst_req_0;
      WPIPE_noblock_obuf_2_2_221_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_2_2_221_inst_req_1;
      WPIPE_noblock_obuf_2_2_221_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_2_219(0);
      data_in <= data_to_outport_205;
      noblock_obuf_2_2_write_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_2_write_1: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_2_2", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_2_2_pipe_write_req(0),
          oack => noblock_obuf_2_2_pipe_write_ack(0),
          odata => noblock_obuf_2_2_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_noblock_obuf_2_3_230_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_2_3_230_inst_req_0;
      WPIPE_noblock_obuf_2_3_230_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_2_3_230_inst_req_1;
      WPIPE_noblock_obuf_2_3_230_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_3_228(0);
      data_in <= data_to_outport_205;
      noblock_obuf_2_3_write_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_3_write_2: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_2_3", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_2_3_pipe_write_req(0),
          oack => noblock_obuf_2_3_pipe_write_ack(0),
          odata => noblock_obuf_2_3_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_noblock_obuf_2_4_239_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_2_4_239_inst_req_0;
      WPIPE_noblock_obuf_2_4_239_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_2_4_239_inst_req_1;
      WPIPE_noblock_obuf_2_4_239_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_4_237(0);
      data_in <= data_to_outport_205;
      noblock_obuf_2_4_write_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_4_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_4_write_3: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_2_4", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_2_4_pipe_write_req(0),
          oack => noblock_obuf_2_4_pipe_write_ack(0),
          odata => noblock_obuf_2_4_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end inputPort_2_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity inputPort_3_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    in_data_3_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_3_pipe_read_data : in   std_logic_vector(31 downto 0);
    noblock_obuf_3_2_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_2_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_3_3_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_3_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_3_4_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_4_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_3_1_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_1_pipe_write_data : out  std_logic_vector(32 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity inputPort_3_Daemon;
architecture inputPort_3_Daemon_arch of inputPort_3_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal inputPort_3_Daemon_CP_407_start: Boolean;
  signal inputPort_3_Daemon_CP_407_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_noblock_obuf_3_2_312_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_3_1_303_inst_req_0 : boolean;
  signal next_count_down_285_254_buf_req_1 : boolean;
  signal WPIPE_noblock_obuf_3_3_321_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_3_2_312_inst_req_1 : boolean;
  signal next_last_dest_id_291_261_buf_ack_0 : boolean;
  signal next_last_dest_id_291_261_buf_ack_1 : boolean;
  signal WPIPE_noblock_obuf_3_3_321_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_3_2_312_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_3_2_312_inst_req_0 : boolean;
  signal next_last_dest_id_291_261_buf_req_1 : boolean;
  signal next_count_down_285_254_buf_ack_0 : boolean;
  signal next_count_down_285_254_buf_req_0 : boolean;
  signal next_last_dest_id_291_261_buf_req_0 : boolean;
  signal phi_stmt_258_req_0 : boolean;
  signal do_while_stmt_248_branch_req_0 : boolean;
  signal WPIPE_noblock_obuf_3_4_330_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_3_4_330_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_3_3_321_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_3_1_303_inst_ack_1 : boolean;
  signal do_while_stmt_248_branch_ack_0 : boolean;
  signal phi_stmt_258_req_1 : boolean;
  signal WPIPE_noblock_obuf_3_3_321_inst_req_1 : boolean;
  signal phi_stmt_250_ack_0 : boolean;
  signal phi_stmt_250_req_0 : boolean;
  signal WPIPE_noblock_obuf_3_1_303_inst_req_1 : boolean;
  signal RPIPE_in_data_3_257_inst_ack_1 : boolean;
  signal RPIPE_in_data_3_257_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_3_4_330_inst_ack_0 : boolean;
  signal RPIPE_in_data_3_257_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_3_4_330_inst_req_0 : boolean;
  signal RPIPE_in_data_3_257_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_3_1_303_inst_ack_0 : boolean;
  signal phi_stmt_258_ack_0 : boolean;
  signal phi_stmt_250_req_1 : boolean;
  signal do_while_stmt_248_branch_ack_1 : boolean;
  signal next_count_down_285_254_buf_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "inputPort_3_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  inputPort_3_Daemon_CP_407_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "inputPort_3_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_3_Daemon_CP_407_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= inputPort_3_Daemon_CP_407_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_3_Daemon_CP_407_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  inputPort_3_Daemon_CP_407: Block -- control-path 
    signal inputPort_3_Daemon_CP_407_elements: BooleanArray(72 downto 0);
    -- 
  begin -- 
    inputPort_3_Daemon_CP_407_elements(0) <= inputPort_3_Daemon_CP_407_start;
    inputPort_3_Daemon_CP_407_symbol <= inputPort_3_Daemon_CP_407_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_247/$entry
      -- CP-element group 0: 	 branch_block_stmt_247/do_while_stmt_248__entry__
      -- CP-element group 0: 	 branch_block_stmt_247/branch_block_stmt_247__entry__
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	72 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_247/$exit
      -- CP-element group 1: 	 branch_block_stmt_247/do_while_stmt_248__exit__
      -- CP-element group 1: 	 branch_block_stmt_247/branch_block_stmt_247__exit__
      -- CP-element group 1: 	 $exit
      -- 
    inputPort_3_Daemon_CP_407_elements(1) <= inputPort_3_Daemon_CP_407_elements(72);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248__entry__
      -- CP-element group 2: 	 branch_block_stmt_247/do_while_stmt_248/$entry
      -- 
    inputPort_3_Daemon_CP_407_elements(2) <= inputPort_3_Daemon_CP_407_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	72 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248__exit__
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_247/do_while_stmt_248/loop_back
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	71 
    -- CP-element group 5: 	70 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_247/do_while_stmt_248/condition_done
      -- CP-element group 5: 	 branch_block_stmt_247/do_while_stmt_248/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_247/do_while_stmt_248/loop_exit/$entry
      -- 
    inputPort_3_Daemon_CP_407_elements(5) <= inputPort_3_Daemon_CP_407_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	69 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_247/do_while_stmt_248/loop_body_done
      -- 
    inputPort_3_Daemon_CP_407_elements(6) <= inputPort_3_Daemon_CP_407_elements(69);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	43 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/back_edge_to_loop_body
      -- 
    inputPort_3_Daemon_CP_407_elements(7) <= inputPort_3_Daemon_CP_407_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	45 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/first_time_through_loop_body
      -- 
    inputPort_3_Daemon_CP_407_elements(8) <= inputPort_3_Daemon_CP_407_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	37 
    -- CP-element group 9: 	38 
    -- CP-element group 9: 	68 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_255_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/$entry
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	68 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/condition_evaluated
      -- 
    condition_evaluated_431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(10), ack => do_while_stmt_248_branch_req_0); -- 
    inputPort_3_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(14) & inputPort_3_Daemon_CP_407_elements(68);
      gj_inputPort_3_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	37 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11: 	39 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_sample_start__ps
      -- 
    inputPort_3_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(9) & inputPort_3_Daemon_CP_407_elements(15) & inputPort_3_Daemon_CP_407_elements(37) & inputPort_3_Daemon_CP_407_elements(14);
      gj_inputPort_3_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	40 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	69 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	37 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_255_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_sample_completed_
      -- 
    inputPort_3_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(17) & inputPort_3_Daemon_CP_407_elements(35) & inputPort_3_Daemon_CP_407_elements(40);
      gj_inputPort_3_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	32 
    -- CP-element group 13: 	38 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13: 	41 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_update_start__ps
      -- 
    inputPort_3_Daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(16) & inputPort_3_Daemon_CP_407_elements(32) & inputPort_3_Daemon_CP_407_elements(38);
      gj_inputPort_3_Daemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	36 
    -- CP-element group 14: 	42 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/aggregated_phi_update_ack
      -- 
    inputPort_3_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(18) & inputPort_3_Daemon_CP_407_elements(36) & inputPort_3_Daemon_CP_407_elements(42);
      gj_inputPort_3_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_sample_start_
      -- 
    inputPort_3_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(9) & inputPort_3_Daemon_CP_407_elements(12);
      gj_inputPort_3_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	57 
    -- CP-element group 16: 	60 
    -- CP-element group 16: 	63 
    -- CP-element group 16: 	66 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_update_start_
      -- 
    inputPort_3_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(9) & inputPort_3_Daemon_CP_407_elements(57) & inputPort_3_Daemon_CP_407_elements(60) & inputPort_3_Daemon_CP_407_elements(63) & inputPort_3_Daemon_CP_407_elements(66);
      gj_inputPort_3_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_sample_completed__ps
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	56 
    -- CP-element group 18: 	59 
    -- CP-element group 18: 	62 
    -- CP-element group 18: 	65 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_update_completed_
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_loopback_trigger
      -- 
    inputPort_3_Daemon_CP_407_elements(19) <= inputPort_3_Daemon_CP_407_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_loopback_sample_req_ps
      -- CP-element group 20: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_loopback_sample_req
      -- 
    phi_stmt_250_loopback_sample_req_446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_250_loopback_sample_req_446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(20), ack => phi_stmt_250_req_1); -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_entry_trigger
      -- 
    inputPort_3_Daemon_CP_407_elements(21) <= inputPort_3_Daemon_CP_407_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_entry_sample_req_ps
      -- CP-element group 22: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_entry_sample_req
      -- 
    phi_stmt_250_entry_sample_req_449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_250_entry_sample_req_449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(22), ack => phi_stmt_250_req_0); -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_phi_mux_ack_ps
      -- CP-element group 23: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_250_phi_mux_ack
      -- 
    phi_stmt_250_phi_mux_ack_452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_250_ack_0, ack => inputPort_3_Daemon_CP_407_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/type_cast_253_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/type_cast_253_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/type_cast_253_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/type_cast_253_sample_start__ps
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/type_cast_253_update_start_
      -- CP-element group 25: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/type_cast_253_update_start__ps
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/type_cast_253_update_completed__ps
      -- 
    inputPort_3_Daemon_CP_407_elements(26) <= inputPort_3_Daemon_CP_407_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/type_cast_253_update_completed_
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => inputPort_3_Daemon_CP_407_elements(25), ack => inputPort_3_Daemon_CP_407_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_Sample/req
      -- CP-element group 28: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_sample_start__ps
      -- 
    req_473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(28), ack => next_count_down_285_254_buf_req_0); -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_Update/req
      -- CP-element group 29: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_update_start_
      -- CP-element group 29: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_update_start__ps
      -- 
    req_478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(29), ack => next_count_down_285_254_buf_req_1); -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_Sample/ack
      -- CP-element group 30: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_sample_completed__ps
      -- 
    ack_474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_285_254_buf_ack_0, ack => inputPort_3_Daemon_CP_407_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_count_down_254_Update/ack
      -- 
    ack_479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_285_254_buf_ack_1, ack => inputPort_3_Daemon_CP_407_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	57 
    -- CP-element group 32: 	60 
    -- CP-element group 32: 	63 
    -- CP-element group 32: 	66 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_255_update_start_
      -- 
    inputPort_3_Daemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(9) & inputPort_3_Daemon_CP_407_elements(57) & inputPort_3_Daemon_CP_407_elements(60) & inputPort_3_Daemon_CP_407_elements(63) & inputPort_3_Daemon_CP_407_elements(66);
      gj_inputPort_3_Daemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/RPIPE_in_data_3_257_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/RPIPE_in_data_3_257_Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/RPIPE_in_data_3_257_Sample/$entry
      -- 
    rr_492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(33), ack => RPIPE_in_data_3_257_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(11) & inputPort_3_Daemon_CP_407_elements(36);
      gj_inputPort_3_Daemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	13 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/RPIPE_in_data_3_257_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/RPIPE_in_data_3_257_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/RPIPE_in_data_3_257_update_start_
      -- 
    cr_497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(34), ack => RPIPE_in_data_3_257_inst_req_1); -- 
    inputPort_3_Daemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(13) & inputPort_3_Daemon_CP_407_elements(35);
      gj_inputPort_3_Daemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/RPIPE_in_data_3_257_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/RPIPE_in_data_3_257_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/RPIPE_in_data_3_257_sample_completed_
      -- 
    ra_493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_3_257_inst_ack_0, ack => inputPort_3_Daemon_CP_407_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	56 
    -- CP-element group 36: 	59 
    -- CP-element group 36: 	62 
    -- CP-element group 36: 	65 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_255_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/RPIPE_in_data_3_257_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/RPIPE_in_data_3_257_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/RPIPE_in_data_3_257_update_completed_
      -- 
    ca_498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_3_257_inst_ack_1, ack => inputPort_3_Daemon_CP_407_elements(36)); -- 
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	9 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	12 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	11 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_sample_start_
      -- 
    inputPort_3_Daemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(9) & inputPort_3_Daemon_CP_407_elements(12);
      gj_inputPort_3_Daemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	9 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	57 
    -- CP-element group 38: 	60 
    -- CP-element group 38: 	63 
    -- CP-element group 38: 	66 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	13 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_update_start_
      -- 
    inputPort_3_Daemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(9) & inputPort_3_Daemon_CP_407_elements(57) & inputPort_3_Daemon_CP_407_elements(60) & inputPort_3_Daemon_CP_407_elements(63) & inputPort_3_Daemon_CP_407_elements(66);
      gj_inputPort_3_Daemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	11 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_sample_start__ps
      -- 
    inputPort_3_Daemon_CP_407_elements(39) <= inputPort_3_Daemon_CP_407_elements(11);
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	12 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_sample_completed__ps
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	13 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_update_start__ps
      -- 
    inputPort_3_Daemon_CP_407_elements(41) <= inputPort_3_Daemon_CP_407_elements(13);
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	14 
    -- CP-element group 42: 	56 
    -- CP-element group 42: 	59 
    -- CP-element group 42: 	62 
    -- CP-element group 42: 	65 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_update_completed__ps
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	7 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_loopback_trigger
      -- 
    inputPort_3_Daemon_CP_407_elements(43) <= inputPort_3_Daemon_CP_407_elements(7);
    -- CP-element group 44:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_loopback_sample_req_ps
      -- CP-element group 44: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_loopback_sample_req
      -- 
    phi_stmt_258_loopback_sample_req_508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_258_loopback_sample_req_508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(44), ack => phi_stmt_258_req_1); -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	8 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_entry_trigger
      -- 
    inputPort_3_Daemon_CP_407_elements(45) <= inputPort_3_Daemon_CP_407_elements(8);
    -- CP-element group 46:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_entry_sample_req_ps
      -- CP-element group 46: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_entry_sample_req
      -- 
    phi_stmt_258_entry_sample_req_511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_258_entry_sample_req_511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(46), ack => phi_stmt_258_req_0); -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_phi_mux_ack_ps
      -- CP-element group 47: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/phi_stmt_258_phi_mux_ack
      -- 
    phi_stmt_258_phi_mux_ack_514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_258_ack_0, ack => inputPort_3_Daemon_CP_407_elements(47)); -- 
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/konst_260_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/konst_260_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/konst_260_sample_completed__ps
      -- CP-element group 48: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/konst_260_sample_start__ps
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/konst_260_update_start__ps
      -- CP-element group 49: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/konst_260_update_start_
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/konst_260_update_completed__ps
      -- 
    inputPort_3_Daemon_CP_407_elements(50) <= inputPort_3_Daemon_CP_407_elements(51);
    -- CP-element group 51:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	50 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/konst_260_update_completed_
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(51) is a control-delay.
    cp_element_51_delay: control_delay_element  generic map(name => " 51_delay", delay_value => 1)  port map(req => inputPort_3_Daemon_CP_407_elements(49), ack => inputPort_3_Daemon_CP_407_elements(51), clk => clk, reset =>reset);
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_Sample/req
      -- CP-element group 52: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_sample_start__ps
      -- 
    req_535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(52), ack => next_last_dest_id_291_261_buf_req_0); -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_Update/req
      -- CP-element group 53: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_update_start_
      -- CP-element group 53: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_update_start__ps
      -- 
    req_540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(53), ack => next_last_dest_id_291_261_buf_req_1); -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_Sample/ack
      -- CP-element group 54: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_sample_completed__ps
      -- 
    ack_536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_291_261_buf_ack_0, ack => inputPort_3_Daemon_CP_407_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_Update/ack
      -- CP-element group 55: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/R_next_last_dest_id_261_update_completed__ps
      -- 
    ack_541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_291_261_buf_ack_1, ack => inputPort_3_Daemon_CP_407_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	18 
    -- CP-element group 56: 	36 
    -- CP-element group 56: 	42 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_1_303_Sample/req
      -- CP-element group 56: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_1_303_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_1_303_sample_start_
      -- 
    req_550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(56), ack => WPIPE_noblock_obuf_3_1_303_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(18) & inputPort_3_Daemon_CP_407_elements(36) & inputPort_3_Daemon_CP_407_elements(42) & inputPort_3_Daemon_CP_407_elements(58);
      gj_inputPort_3_Daemon_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	16 
    -- CP-element group 57: 	32 
    -- CP-element group 57: 	38 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_1_303_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_1_303_update_start_
      -- CP-element group 57: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_1_303_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_1_303_Update/req
      -- CP-element group 57: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_1_303_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_1_303_Sample/ack
      -- 
    ack_551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_1_303_inst_ack_0, ack => inputPort_3_Daemon_CP_407_elements(57)); -- 
    req_555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(57), ack => WPIPE_noblock_obuf_3_1_303_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	69 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_1_303_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_1_303_Update/ack
      -- CP-element group 58: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_1_303_Update/$exit
      -- 
    ack_556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_1_303_inst_ack_1, ack => inputPort_3_Daemon_CP_407_elements(58)); -- 
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	18 
    -- CP-element group 59: 	36 
    -- CP-element group 59: 	42 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_2_312_Sample/req
      -- CP-element group 59: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_2_312_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_2_312_sample_start_
      -- 
    req_564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(59), ack => WPIPE_noblock_obuf_3_2_312_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(18) & inputPort_3_Daemon_CP_407_elements(36) & inputPort_3_Daemon_CP_407_elements(42) & inputPort_3_Daemon_CP_407_elements(61);
      gj_inputPort_3_Daemon_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	16 
    -- CP-element group 60: 	32 
    -- CP-element group 60: 	38 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_2_312_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_2_312_Update/req
      -- CP-element group 60: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_2_312_Sample/ack
      -- CP-element group 60: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_2_312_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_2_312_update_start_
      -- CP-element group 60: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_2_312_sample_completed_
      -- 
    ack_565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_2_312_inst_ack_0, ack => inputPort_3_Daemon_CP_407_elements(60)); -- 
    req_569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(60), ack => WPIPE_noblock_obuf_3_2_312_inst_req_1); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	69 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_2_312_Update/ack
      -- CP-element group 61: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_2_312_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_2_312_update_completed_
      -- 
    ack_570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_2_312_inst_ack_1, ack => inputPort_3_Daemon_CP_407_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	18 
    -- CP-element group 62: 	36 
    -- CP-element group 62: 	42 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_3_321_Sample/req
      -- CP-element group 62: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_3_321_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_3_321_sample_start_
      -- 
    req_578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(62), ack => WPIPE_noblock_obuf_3_3_321_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(18) & inputPort_3_Daemon_CP_407_elements(36) & inputPort_3_Daemon_CP_407_elements(42) & inputPort_3_Daemon_CP_407_elements(64);
      gj_inputPort_3_Daemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	16 
    -- CP-element group 63: 	32 
    -- CP-element group 63: 	38 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_3_321_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_3_321_Sample/ack
      -- CP-element group 63: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_3_321_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_3_321_Update/req
      -- CP-element group 63: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_3_321_update_start_
      -- CP-element group 63: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_3_321_sample_completed_
      -- 
    ack_579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_3_321_inst_ack_0, ack => inputPort_3_Daemon_CP_407_elements(63)); -- 
    req_583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(63), ack => WPIPE_noblock_obuf_3_3_321_inst_req_1); -- 
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	69 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_3_321_Update/ack
      -- CP-element group 64: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_3_321_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_3_321_Update/$exit
      -- 
    ack_584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_3_321_inst_ack_1, ack => inputPort_3_Daemon_CP_407_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	18 
    -- CP-element group 65: 	36 
    -- CP-element group 65: 	42 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_4_330_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_4_330_Sample/req
      -- CP-element group 65: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_4_330_Sample/$entry
      -- 
    req_592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(65), ack => WPIPE_noblock_obuf_3_4_330_inst_req_0); -- 
    inputPort_3_Daemon_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(18) & inputPort_3_Daemon_CP_407_elements(36) & inputPort_3_Daemon_CP_407_elements(42) & inputPort_3_Daemon_CP_407_elements(67);
      gj_inputPort_3_Daemon_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	16 
    -- CP-element group 66: 	32 
    -- CP-element group 66: 	38 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_4_330_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_4_330_update_start_
      -- CP-element group 66: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_4_330_Update/req
      -- CP-element group 66: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_4_330_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_4_330_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_4_330_Sample/$exit
      -- 
    ack_593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_4_330_inst_ack_0, ack => inputPort_3_Daemon_CP_407_elements(66)); -- 
    req_597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_3_Daemon_CP_407_elements(66), ack => WPIPE_noblock_obuf_3_4_330_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_4_330_Update/ack
      -- CP-element group 67: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_4_330_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/WPIPE_noblock_obuf_3_4_330_Update/$exit
      -- 
    ack_598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_3_4_330_inst_ack_1, ack => inputPort_3_Daemon_CP_407_elements(67)); -- 
    -- CP-element group 68:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	9 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	10 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group inputPort_3_Daemon_CP_407_elements(68) is a control-delay.
    cp_element_68_delay: control_delay_element  generic map(name => " 68_delay", delay_value => 1)  port map(req => inputPort_3_Daemon_CP_407_elements(9), ack => inputPort_3_Daemon_CP_407_elements(68), clk => clk, reset =>reset);
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	12 
    -- CP-element group 69: 	58 
    -- CP-element group 69: 	61 
    -- CP-element group 69: 	64 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	6 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_247/do_while_stmt_248/do_while_stmt_248_loop_body/$exit
      -- 
    inputPort_3_Daemon_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_3_Daemon_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_3_Daemon_CP_407_elements(12) & inputPort_3_Daemon_CP_407_elements(58) & inputPort_3_Daemon_CP_407_elements(61) & inputPort_3_Daemon_CP_407_elements(64) & inputPort_3_Daemon_CP_407_elements(67);
      gj_inputPort_3_Daemon_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	5 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_247/do_while_stmt_248/loop_exit/ack
      -- CP-element group 70: 	 branch_block_stmt_247/do_while_stmt_248/loop_exit/$exit
      -- 
    ack_603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_248_branch_ack_0, ack => inputPort_3_Daemon_CP_407_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	5 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_247/do_while_stmt_248/loop_taken/$exit
      -- CP-element group 71: 	 branch_block_stmt_247/do_while_stmt_248/loop_taken/ack
      -- 
    ack_607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_248_branch_ack_1, ack => inputPort_3_Daemon_CP_407_elements(71)); -- 
    -- CP-element group 72:  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	3 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	1 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_247/do_while_stmt_248/$exit
      -- 
    inputPort_3_Daemon_CP_407_elements(72) <= inputPort_3_Daemon_CP_407_elements(3);
    inputPort_3_Daemon_do_while_stmt_248_terminator_608: loop_terminator -- 
      generic map (name => " inputPort_3_Daemon_do_while_stmt_248_terminator_608", max_iterations_in_flight =>7) 
      port map(loop_body_exit => inputPort_3_Daemon_CP_407_elements(6),loop_continue => inputPort_3_Daemon_CP_407_elements(71),loop_terminate => inputPort_3_Daemon_CP_407_elements(70),loop_back => inputPort_3_Daemon_CP_407_elements(4),loop_exit => inputPort_3_Daemon_CP_407_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_250_phi_seq_480_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_3_Daemon_CP_407_elements(21);
      inputPort_3_Daemon_CP_407_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_3_Daemon_CP_407_elements(24);
      inputPort_3_Daemon_CP_407_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_3_Daemon_CP_407_elements(26);
      inputPort_3_Daemon_CP_407_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_3_Daemon_CP_407_elements(19);
      inputPort_3_Daemon_CP_407_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_3_Daemon_CP_407_elements(30);
      inputPort_3_Daemon_CP_407_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_3_Daemon_CP_407_elements(31);
      inputPort_3_Daemon_CP_407_elements(20) <= phi_mux_reqs(1);
      phi_stmt_250_phi_seq_480 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_250_phi_seq_480") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_3_Daemon_CP_407_elements(11), 
          phi_sample_ack => inputPort_3_Daemon_CP_407_elements(17), 
          phi_update_req => inputPort_3_Daemon_CP_407_elements(13), 
          phi_update_ack => inputPort_3_Daemon_CP_407_elements(18), 
          phi_mux_ack => inputPort_3_Daemon_CP_407_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_258_phi_seq_542_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_3_Daemon_CP_407_elements(45);
      inputPort_3_Daemon_CP_407_elements(48)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_3_Daemon_CP_407_elements(48);
      inputPort_3_Daemon_CP_407_elements(49)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_3_Daemon_CP_407_elements(50);
      inputPort_3_Daemon_CP_407_elements(46) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_3_Daemon_CP_407_elements(43);
      inputPort_3_Daemon_CP_407_elements(52)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_3_Daemon_CP_407_elements(54);
      inputPort_3_Daemon_CP_407_elements(53)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_3_Daemon_CP_407_elements(55);
      inputPort_3_Daemon_CP_407_elements(44) <= phi_mux_reqs(1);
      phi_stmt_258_phi_seq_542 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_258_phi_seq_542") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_3_Daemon_CP_407_elements(39), 
          phi_sample_ack => inputPort_3_Daemon_CP_407_elements(40), 
          phi_update_req => inputPort_3_Daemon_CP_407_elements(41), 
          phi_update_ack => inputPort_3_Daemon_CP_407_elements(42), 
          phi_mux_ack => inputPort_3_Daemon_CP_407_elements(47), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_432_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= inputPort_3_Daemon_CP_407_elements(7);
        preds(1)  <= inputPort_3_Daemon_CP_407_elements(8);
        entry_tmerge_432 : transition_merge -- 
          generic map(name => " entry_tmerge_432")
          port map (preds => preds, symbol_out => inputPort_3_Daemon_CP_407_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal RPIPE_in_data_3_257_wire : std_logic_vector(31 downto 0);
    signal R_ONE_1_293_wire_constant : std_logic_vector(0 downto 0);
    signal SUB_u16_u16_280_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_283_wire : std_logic_vector(15 downto 0);
    signal count_down_250 : std_logic_vector(15 downto 0);
    signal data_to_outport_296 : std_logic_vector(32 downto 0);
    signal dest_id_271 : std_logic_vector(7 downto 0);
    signal input_word_255 : std_logic_vector(31 downto 0);
    signal konst_260_wire_constant : std_logic_vector(7 downto 0);
    signal konst_265_wire_constant : std_logic_vector(15 downto 0);
    signal konst_279_wire_constant : std_logic_vector(15 downto 0);
    signal konst_282_wire_constant : std_logic_vector(15 downto 0);
    signal konst_299_wire_constant : std_logic_vector(7 downto 0);
    signal konst_308_wire_constant : std_logic_vector(7 downto 0);
    signal konst_317_wire_constant : std_logic_vector(7 downto 0);
    signal konst_326_wire_constant : std_logic_vector(7 downto 0);
    signal konst_334_wire_constant : std_logic_vector(0 downto 0);
    signal last_dest_id_258 : std_logic_vector(7 downto 0);
    signal new_packet_267 : std_logic_vector(0 downto 0);
    signal next_count_down_285 : std_logic_vector(15 downto 0);
    signal next_count_down_285_254_buffered : std_logic_vector(15 downto 0);
    signal next_last_dest_id_291 : std_logic_vector(7 downto 0);
    signal next_last_dest_id_291_261_buffered : std_logic_vector(7 downto 0);
    signal pkt_length_275 : std_logic_vector(15 downto 0);
    signal send_to_1_301 : std_logic_vector(0 downto 0);
    signal send_to_2_310 : std_logic_vector(0 downto 0);
    signal send_to_3_319 : std_logic_vector(0 downto 0);
    signal send_to_4_328 : std_logic_vector(0 downto 0);
    signal type_cast_253_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    R_ONE_1_293_wire_constant <= "1";
    konst_260_wire_constant <= "00000000";
    konst_265_wire_constant <= "0000000000000000";
    konst_279_wire_constant <= "0000000000000001";
    konst_282_wire_constant <= "0000000000000001";
    konst_299_wire_constant <= "00000001";
    konst_308_wire_constant <= "00000010";
    konst_317_wire_constant <= "00000011";
    konst_326_wire_constant <= "00000100";
    konst_334_wire_constant <= "1";
    type_cast_253_wire_constant <= "0000000000000000";
    phi_stmt_250: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_253_wire_constant & next_count_down_285_254_buffered;
      req <= phi_stmt_250_req_0 & phi_stmt_250_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_250",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_250_ack_0,
          idata => idata,
          odata => count_down_250,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_250
    phi_stmt_258: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_260_wire_constant & next_last_dest_id_291_261_buffered;
      req <= phi_stmt_258_req_0 & phi_stmt_258_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_258",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_258_ack_0,
          idata => idata,
          odata => last_dest_id_258,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_258
    -- flow-through select operator MUX_284_inst
    next_count_down_285 <= SUB_u16_u16_280_wire when (new_packet_267(0) /=  '0') else SUB_u16_u16_283_wire;
    -- flow-through select operator MUX_290_inst
    next_last_dest_id_291 <= dest_id_271 when (new_packet_267(0) /=  '0') else last_dest_id_258;
    -- flow-through slice operator slice_270_inst
    dest_id_271 <= input_word_255(31 downto 24);
    -- flow-through slice operator slice_274_inst
    pkt_length_275 <= input_word_255(23 downto 8);
    next_count_down_285_254_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_count_down_285_254_buf_req_0;
      next_count_down_285_254_buf_ack_0<= wack(0);
      rreq(0) <= next_count_down_285_254_buf_req_1;
      next_count_down_285_254_buf_ack_1<= rack(0);
      next_count_down_285_254_buf : InterlockBuffer generic map ( -- 
        name => "next_count_down_285_254_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_count_down_285,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_count_down_285_254_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_last_dest_id_291_261_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_last_dest_id_291_261_buf_req_0;
      next_last_dest_id_291_261_buf_ack_0<= wack(0);
      rreq(0) <= next_last_dest_id_291_261_buf_req_1;
      next_last_dest_id_291_261_buf_ack_1<= rack(0);
      next_last_dest_id_291_261_buf : InterlockBuffer generic map ( -- 
        name => "next_last_dest_id_291_261_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_last_dest_id_291,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_last_dest_id_291_261_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_255
    process(RPIPE_in_data_3_257_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := RPIPE_in_data_3_257_wire(31 downto 0);
      input_word_255 <= tmp_var; -- 
    end process;
    do_while_stmt_248_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_334_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_248_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_248_branch_req_0,
          ack0 => do_while_stmt_248_branch_ack_0,
          ack1 => do_while_stmt_248_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator CONCAT_u1_u33_295_inst
    process(R_ONE_1_293_wire_constant, input_word_255) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ONE_1_293_wire_constant, input_word_255, tmp_var);
      data_to_outport_296 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_266_inst
    process(count_down_250) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(count_down_250, konst_265_wire_constant, tmp_var);
      new_packet_267 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_300_inst
    process(next_last_dest_id_291) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_291, konst_299_wire_constant, tmp_var);
      send_to_1_301 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_309_inst
    process(next_last_dest_id_291) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_291, konst_308_wire_constant, tmp_var);
      send_to_2_310 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_318_inst
    process(next_last_dest_id_291) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_291, konst_317_wire_constant, tmp_var);
      send_to_3_319 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_327_inst
    process(next_last_dest_id_291) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_291, konst_326_wire_constant, tmp_var);
      send_to_4_328 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_280_inst
    process(pkt_length_275) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(pkt_length_275, konst_279_wire_constant, tmp_var);
      SUB_u16_u16_280_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_283_inst
    process(count_down_250) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(count_down_250, konst_282_wire_constant, tmp_var);
      SUB_u16_u16_283_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_in_data_3_257_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_in_data_3_257_inst_req_0;
      RPIPE_in_data_3_257_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_in_data_3_257_inst_req_1;
      RPIPE_in_data_3_257_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_in_data_3_257_wire <= data_out(31 downto 0);
      in_data_3_read_0_gI: SplitGuardInterface generic map(name => "in_data_3_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      in_data_3_read_0: InputPortRevised -- 
        generic map ( name => "in_data_3_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => in_data_3_pipe_read_req(0),
          oack => in_data_3_pipe_read_ack(0),
          odata => in_data_3_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_noblock_obuf_3_1_303_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_3_1_303_inst_req_0;
      WPIPE_noblock_obuf_3_1_303_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_3_1_303_inst_req_1;
      WPIPE_noblock_obuf_3_1_303_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_1_301(0);
      data_in <= data_to_outport_296;
      noblock_obuf_3_1_write_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_1_write_0: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_3_1", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_3_1_pipe_write_req(0),
          oack => noblock_obuf_3_1_pipe_write_ack(0),
          odata => noblock_obuf_3_1_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_noblock_obuf_3_2_312_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_3_2_312_inst_req_0;
      WPIPE_noblock_obuf_3_2_312_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_3_2_312_inst_req_1;
      WPIPE_noblock_obuf_3_2_312_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_2_310(0);
      data_in <= data_to_outport_296;
      noblock_obuf_3_2_write_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_2_write_1: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_3_2", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_3_2_pipe_write_req(0),
          oack => noblock_obuf_3_2_pipe_write_ack(0),
          odata => noblock_obuf_3_2_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_noblock_obuf_3_3_321_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_3_3_321_inst_req_0;
      WPIPE_noblock_obuf_3_3_321_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_3_3_321_inst_req_1;
      WPIPE_noblock_obuf_3_3_321_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_3_319(0);
      data_in <= data_to_outport_296;
      noblock_obuf_3_3_write_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_3_write_2: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_3_3", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_3_3_pipe_write_req(0),
          oack => noblock_obuf_3_3_pipe_write_ack(0),
          odata => noblock_obuf_3_3_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_noblock_obuf_3_4_330_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_3_4_330_inst_req_0;
      WPIPE_noblock_obuf_3_4_330_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_3_4_330_inst_req_1;
      WPIPE_noblock_obuf_3_4_330_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_4_328(0);
      data_in <= data_to_outport_296;
      noblock_obuf_3_4_write_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_4_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_4_write_3: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_3_4", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_3_4_pipe_write_req(0),
          oack => noblock_obuf_3_4_pipe_write_ack(0),
          odata => noblock_obuf_3_4_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end inputPort_3_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity inputPort_4_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    in_data_4_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_4_pipe_read_data : in   std_logic_vector(31 downto 0);
    noblock_obuf_4_1_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_1_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_4_2_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_2_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_4_3_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_3_pipe_write_data : out  std_logic_vector(32 downto 0);
    noblock_obuf_4_4_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_4_pipe_write_data : out  std_logic_vector(32 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity inputPort_4_Daemon;
architecture inputPort_4_Daemon_arch of inputPort_4_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal inputPort_4_Daemon_CP_609_start: Boolean;
  signal inputPort_4_Daemon_CP_609_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_339_branch_req_0 : boolean;
  signal phi_stmt_341_req_1 : boolean;
  signal phi_stmt_341_req_0 : boolean;
  signal phi_stmt_341_ack_0 : boolean;
  signal next_count_down_376_345_buf_req_0 : boolean;
  signal next_count_down_376_345_buf_ack_0 : boolean;
  signal next_count_down_376_345_buf_req_1 : boolean;
  signal next_count_down_376_345_buf_ack_1 : boolean;
  signal RPIPE_in_data_4_348_inst_req_0 : boolean;
  signal RPIPE_in_data_4_348_inst_ack_0 : boolean;
  signal RPIPE_in_data_4_348_inst_req_1 : boolean;
  signal RPIPE_in_data_4_348_inst_ack_1 : boolean;
  signal phi_stmt_349_req_1 : boolean;
  signal phi_stmt_349_req_0 : boolean;
  signal phi_stmt_349_ack_0 : boolean;
  signal next_last_dest_id_382_352_buf_req_0 : boolean;
  signal next_last_dest_id_382_352_buf_ack_0 : boolean;
  signal next_last_dest_id_382_352_buf_req_1 : boolean;
  signal next_last_dest_id_382_352_buf_ack_1 : boolean;
  signal WPIPE_noblock_obuf_4_1_394_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_4_1_394_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_4_1_394_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_4_1_394_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_4_2_403_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_4_2_403_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_4_2_403_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_4_2_403_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_4_3_412_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_4_3_412_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_4_3_412_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_4_3_412_inst_ack_1 : boolean;
  signal WPIPE_noblock_obuf_4_4_421_inst_req_0 : boolean;
  signal WPIPE_noblock_obuf_4_4_421_inst_ack_0 : boolean;
  signal WPIPE_noblock_obuf_4_4_421_inst_req_1 : boolean;
  signal WPIPE_noblock_obuf_4_4_421_inst_ack_1 : boolean;
  signal do_while_stmt_339_branch_ack_0 : boolean;
  signal do_while_stmt_339_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "inputPort_4_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  inputPort_4_Daemon_CP_609_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "inputPort_4_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_4_Daemon_CP_609_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= inputPort_4_Daemon_CP_609_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= inputPort_4_Daemon_CP_609_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  inputPort_4_Daemon_CP_609: Block -- control-path 
    signal inputPort_4_Daemon_CP_609_elements: BooleanArray(72 downto 0);
    -- 
  begin -- 
    inputPort_4_Daemon_CP_609_elements(0) <= inputPort_4_Daemon_CP_609_start;
    inputPort_4_Daemon_CP_609_symbol <= inputPort_4_Daemon_CP_609_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_338/branch_block_stmt_338__entry__
      -- CP-element group 0: 	 branch_block_stmt_338/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_338/do_while_stmt_339__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	72 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_338/branch_block_stmt_338__exit__
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_338/$exit
      -- CP-element group 1: 	 branch_block_stmt_338/do_while_stmt_339__exit__
      -- 
    inputPort_4_Daemon_CP_609_elements(1) <= inputPort_4_Daemon_CP_609_elements(72);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339__entry__
      -- CP-element group 2: 	 branch_block_stmt_338/do_while_stmt_339/$entry
      -- 
    inputPort_4_Daemon_CP_609_elements(2) <= inputPort_4_Daemon_CP_609_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	72 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339__exit__
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_338/do_while_stmt_339/loop_back
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	71 
    -- CP-element group 5: 	70 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_338/do_while_stmt_339/condition_done
      -- CP-element group 5: 	 branch_block_stmt_338/do_while_stmt_339/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_338/do_while_stmt_339/loop_taken/$entry
      -- 
    inputPort_4_Daemon_CP_609_elements(5) <= inputPort_4_Daemon_CP_609_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	69 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_338/do_while_stmt_339/loop_body_done
      -- 
    inputPort_4_Daemon_CP_609_elements(6) <= inputPort_4_Daemon_CP_609_elements(69);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	43 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/back_edge_to_loop_body
      -- 
    inputPort_4_Daemon_CP_609_elements(7) <= inputPort_4_Daemon_CP_609_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	45 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/first_time_through_loop_body
      -- 
    inputPort_4_Daemon_CP_609_elements(8) <= inputPort_4_Daemon_CP_609_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	68 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	37 
    -- CP-element group 9: 	38 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_346_sample_start_
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	68 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/condition_evaluated
      -- 
    condition_evaluated_633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(10), ack => do_while_stmt_339_branch_req_0); -- 
    inputPort_4_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(68) & inputPort_4_Daemon_CP_609_elements(14);
      gj_inputPort_4_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	37 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11: 	39 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_sample_start__ps
      -- 
    inputPort_4_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(9) & inputPort_4_Daemon_CP_609_elements(15) & inputPort_4_Daemon_CP_609_elements(37) & inputPort_4_Daemon_CP_609_elements(14);
      gj_inputPort_4_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	40 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	69 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	37 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_346_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_sample_completed_
      -- 
    inputPort_4_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(17) & inputPort_4_Daemon_CP_609_elements(35) & inputPort_4_Daemon_CP_609_elements(40);
      gj_inputPort_4_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	32 
    -- CP-element group 13: 	38 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13: 	41 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/aggregated_phi_update_req
      -- 
    inputPort_4_Daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(16) & inputPort_4_Daemon_CP_609_elements(32) & inputPort_4_Daemon_CP_609_elements(38);
      gj_inputPort_4_Daemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	36 
    -- CP-element group 14: 	42 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/aggregated_phi_update_ack
      -- 
    inputPort_4_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(18) & inputPort_4_Daemon_CP_609_elements(36) & inputPort_4_Daemon_CP_609_elements(42);
      gj_inputPort_4_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_sample_start_
      -- 
    inputPort_4_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(9) & inputPort_4_Daemon_CP_609_elements(12);
      gj_inputPort_4_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	66 
    -- CP-element group 16: 	60 
    -- CP-element group 16: 	63 
    -- CP-element group 16: 	57 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_update_start_
      -- 
    inputPort_4_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(9) & inputPort_4_Daemon_CP_609_elements(66) & inputPort_4_Daemon_CP_609_elements(60) & inputPort_4_Daemon_CP_609_elements(63) & inputPort_4_Daemon_CP_609_elements(57);
      gj_inputPort_4_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_sample_completed__ps
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	56 
    -- CP-element group 18: 	59 
    -- CP-element group 18: 	65 
    -- CP-element group 18: 	62 
    -- CP-element group 18: 	14 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_update_completed_
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_loopback_trigger
      -- 
    inputPort_4_Daemon_CP_609_elements(19) <= inputPort_4_Daemon_CP_609_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_loopback_sample_req_ps
      -- 
    phi_stmt_341_loopback_sample_req_648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_341_loopback_sample_req_648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(20), ack => phi_stmt_341_req_1); -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_entry_trigger
      -- 
    inputPort_4_Daemon_CP_609_elements(21) <= inputPort_4_Daemon_CP_609_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_entry_sample_req_ps
      -- 
    phi_stmt_341_entry_sample_req_651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_341_entry_sample_req_651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(22), ack => phi_stmt_341_req_0); -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_341_phi_mux_ack_ps
      -- 
    phi_stmt_341_phi_mux_ack_654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_341_ack_0, ack => inputPort_4_Daemon_CP_609_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/type_cast_344_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/type_cast_344_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/type_cast_344_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/type_cast_344_sample_completed_
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/type_cast_344_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/type_cast_344_update_start_
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/type_cast_344_update_completed__ps
      -- 
    inputPort_4_Daemon_CP_609_elements(26) <= inputPort_4_Daemon_CP_609_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/type_cast_344_update_completed_
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => inputPort_4_Daemon_CP_609_elements(25), ack => inputPort_4_Daemon_CP_609_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_Sample/req
      -- 
    req_675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(28), ack => next_count_down_376_345_buf_req_0); -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_update_start_
      -- CP-element group 29: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_Update/req
      -- 
    req_680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(29), ack => next_count_down_376_345_buf_req_1); -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_Sample/ack
      -- 
    ack_676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_376_345_buf_ack_0, ack => inputPort_4_Daemon_CP_609_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_count_down_345_Update/ack
      -- 
    ack_681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_down_376_345_buf_ack_1, ack => inputPort_4_Daemon_CP_609_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	66 
    -- CP-element group 32: 	60 
    -- CP-element group 32: 	63 
    -- CP-element group 32: 	57 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_346_update_start_
      -- 
    inputPort_4_Daemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(9) & inputPort_4_Daemon_CP_609_elements(66) & inputPort_4_Daemon_CP_609_elements(60) & inputPort_4_Daemon_CP_609_elements(63) & inputPort_4_Daemon_CP_609_elements(57);
      gj_inputPort_4_Daemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/RPIPE_in_data_4_348_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/RPIPE_in_data_4_348_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/RPIPE_in_data_4_348_Sample/rr
      -- 
    rr_694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(33), ack => RPIPE_in_data_4_348_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(11) & inputPort_4_Daemon_CP_609_elements(36);
      gj_inputPort_4_Daemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	13 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/RPIPE_in_data_4_348_update_start_
      -- CP-element group 34: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/RPIPE_in_data_4_348_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/RPIPE_in_data_4_348_Update/cr
      -- 
    cr_699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(34), ack => RPIPE_in_data_4_348_inst_req_1); -- 
    inputPort_4_Daemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(13) & inputPort_4_Daemon_CP_609_elements(35);
      gj_inputPort_4_Daemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/RPIPE_in_data_4_348_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/RPIPE_in_data_4_348_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/RPIPE_in_data_4_348_Sample/ra
      -- 
    ra_695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_4_348_inst_ack_0, ack => inputPort_4_Daemon_CP_609_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	56 
    -- CP-element group 36: 	59 
    -- CP-element group 36: 	65 
    -- CP-element group 36: 	62 
    -- CP-element group 36: 	14 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_346_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/RPIPE_in_data_4_348_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/RPIPE_in_data_4_348_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/RPIPE_in_data_4_348_Update/ca
      -- 
    ca_700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_in_data_4_348_inst_ack_1, ack => inputPort_4_Daemon_CP_609_elements(36)); -- 
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	9 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	12 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	11 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_sample_start_
      -- 
    inputPort_4_Daemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(9) & inputPort_4_Daemon_CP_609_elements(12);
      gj_inputPort_4_Daemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	9 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	66 
    -- CP-element group 38: 	60 
    -- CP-element group 38: 	63 
    -- CP-element group 38: 	57 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	13 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_update_start_
      -- 
    inputPort_4_Daemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(9) & inputPort_4_Daemon_CP_609_elements(66) & inputPort_4_Daemon_CP_609_elements(60) & inputPort_4_Daemon_CP_609_elements(63) & inputPort_4_Daemon_CP_609_elements(57);
      gj_inputPort_4_Daemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	11 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_sample_start__ps
      -- 
    inputPort_4_Daemon_CP_609_elements(39) <= inputPort_4_Daemon_CP_609_elements(11);
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	12 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_sample_completed__ps
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	13 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_update_start__ps
      -- 
    inputPort_4_Daemon_CP_609_elements(41) <= inputPort_4_Daemon_CP_609_elements(13);
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	56 
    -- CP-element group 42: 	59 
    -- CP-element group 42: 	65 
    -- CP-element group 42: 	62 
    -- CP-element group 42: 	14 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_update_completed__ps
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	7 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_loopback_trigger
      -- 
    inputPort_4_Daemon_CP_609_elements(43) <= inputPort_4_Daemon_CP_609_elements(7);
    -- CP-element group 44:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_loopback_sample_req
      -- CP-element group 44: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_loopback_sample_req_ps
      -- 
    phi_stmt_349_loopback_sample_req_710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_349_loopback_sample_req_710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(44), ack => phi_stmt_349_req_1); -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	8 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_entry_trigger
      -- 
    inputPort_4_Daemon_CP_609_elements(45) <= inputPort_4_Daemon_CP_609_elements(8);
    -- CP-element group 46:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_entry_sample_req
      -- CP-element group 46: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_entry_sample_req_ps
      -- 
    phi_stmt_349_entry_sample_req_713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_349_entry_sample_req_713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(46), ack => phi_stmt_349_req_0); -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_phi_mux_ack
      -- CP-element group 47: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/phi_stmt_349_phi_mux_ack_ps
      -- 
    phi_stmt_349_phi_mux_ack_716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_349_ack_0, ack => inputPort_4_Daemon_CP_609_elements(47)); -- 
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/konst_351_sample_start__ps
      -- CP-element group 48: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/konst_351_sample_completed__ps
      -- CP-element group 48: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/konst_351_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/konst_351_sample_completed_
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/konst_351_update_start__ps
      -- CP-element group 49: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/konst_351_update_start_
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/konst_351_update_completed__ps
      -- 
    inputPort_4_Daemon_CP_609_elements(50) <= inputPort_4_Daemon_CP_609_elements(51);
    -- CP-element group 51:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	50 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/konst_351_update_completed_
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(51) is a control-delay.
    cp_element_51_delay: control_delay_element  generic map(name => " 51_delay", delay_value => 1)  port map(req => inputPort_4_Daemon_CP_609_elements(49), ack => inputPort_4_Daemon_CP_609_elements(51), clk => clk, reset =>reset);
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_Sample/req
      -- 
    req_737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(52), ack => next_last_dest_id_382_352_buf_req_0); -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_update_start_
      -- CP-element group 53: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_Update/req
      -- 
    req_742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(53), ack => next_last_dest_id_382_352_buf_req_1); -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_Sample/ack
      -- 
    ack_738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_382_352_buf_ack_0, ack => inputPort_4_Daemon_CP_609_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/R_next_last_dest_id_352_Update/ack
      -- 
    ack_743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_last_dest_id_382_352_buf_ack_1, ack => inputPort_4_Daemon_CP_609_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	18 
    -- CP-element group 56: 	36 
    -- CP-element group 56: 	42 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_1_394_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_1_394_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_1_394_Sample/req
      -- 
    req_752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(56), ack => WPIPE_noblock_obuf_4_1_394_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(18) & inputPort_4_Daemon_CP_609_elements(36) & inputPort_4_Daemon_CP_609_elements(42) & inputPort_4_Daemon_CP_609_elements(58);
      gj_inputPort_4_Daemon_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	16 
    -- CP-element group 57: 	32 
    -- CP-element group 57: 	38 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_1_394_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_1_394_update_start_
      -- CP-element group 57: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_1_394_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_1_394_Sample/ack
      -- CP-element group 57: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_1_394_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_1_394_Update/req
      -- 
    ack_753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_1_394_inst_ack_0, ack => inputPort_4_Daemon_CP_609_elements(57)); -- 
    req_757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(57), ack => WPIPE_noblock_obuf_4_1_394_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	69 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_1_394_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_1_394_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_1_394_Update/ack
      -- 
    ack_758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_1_394_inst_ack_1, ack => inputPort_4_Daemon_CP_609_elements(58)); -- 
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	18 
    -- CP-element group 59: 	36 
    -- CP-element group 59: 	42 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_2_403_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_2_403_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_2_403_Sample/req
      -- 
    req_766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(59), ack => WPIPE_noblock_obuf_4_2_403_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(18) & inputPort_4_Daemon_CP_609_elements(36) & inputPort_4_Daemon_CP_609_elements(42) & inputPort_4_Daemon_CP_609_elements(61);
      gj_inputPort_4_Daemon_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	16 
    -- CP-element group 60: 	32 
    -- CP-element group 60: 	38 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_2_403_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_2_403_update_start_
      -- CP-element group 60: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_2_403_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_2_403_Sample/ack
      -- CP-element group 60: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_2_403_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_2_403_Update/req
      -- 
    ack_767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_2_403_inst_ack_0, ack => inputPort_4_Daemon_CP_609_elements(60)); -- 
    req_771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(60), ack => WPIPE_noblock_obuf_4_2_403_inst_req_1); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	69 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_2_403_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_2_403_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_2_403_Update/ack
      -- 
    ack_772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_2_403_inst_ack_1, ack => inputPort_4_Daemon_CP_609_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	18 
    -- CP-element group 62: 	36 
    -- CP-element group 62: 	42 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_3_412_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_3_412_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_3_412_Sample/req
      -- 
    req_780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(62), ack => WPIPE_noblock_obuf_4_3_412_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(18) & inputPort_4_Daemon_CP_609_elements(36) & inputPort_4_Daemon_CP_609_elements(42) & inputPort_4_Daemon_CP_609_elements(64);
      gj_inputPort_4_Daemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	16 
    -- CP-element group 63: 	32 
    -- CP-element group 63: 	38 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_3_412_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_3_412_update_start_
      -- CP-element group 63: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_3_412_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_3_412_Sample/ack
      -- CP-element group 63: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_3_412_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_3_412_Update/req
      -- 
    ack_781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_3_412_inst_ack_0, ack => inputPort_4_Daemon_CP_609_elements(63)); -- 
    req_785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(63), ack => WPIPE_noblock_obuf_4_3_412_inst_req_1); -- 
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	69 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_3_412_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_3_412_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_3_412_Update/ack
      -- 
    ack_786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_3_412_inst_ack_1, ack => inputPort_4_Daemon_CP_609_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	18 
    -- CP-element group 65: 	36 
    -- CP-element group 65: 	42 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_4_421_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_4_421_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_4_421_Sample/req
      -- 
    req_794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(65), ack => WPIPE_noblock_obuf_4_4_421_inst_req_0); -- 
    inputPort_4_Daemon_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(18) & inputPort_4_Daemon_CP_609_elements(36) & inputPort_4_Daemon_CP_609_elements(42) & inputPort_4_Daemon_CP_609_elements(67);
      gj_inputPort_4_Daemon_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	16 
    -- CP-element group 66: 	32 
    -- CP-element group 66: 	38 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_4_421_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_4_421_update_start_
      -- CP-element group 66: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_4_421_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_4_421_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_4_421_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_4_421_Update/req
      -- 
    ack_795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_4_421_inst_ack_0, ack => inputPort_4_Daemon_CP_609_elements(66)); -- 
    req_799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => inputPort_4_Daemon_CP_609_elements(66), ack => WPIPE_noblock_obuf_4_4_421_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_4_421_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_4_421_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/WPIPE_noblock_obuf_4_4_421_Update/ack
      -- 
    ack_800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_noblock_obuf_4_4_421_inst_ack_1, ack => inputPort_4_Daemon_CP_609_elements(67)); -- 
    -- CP-element group 68:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	9 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	10 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group inputPort_4_Daemon_CP_609_elements(68) is a control-delay.
    cp_element_68_delay: control_delay_element  generic map(name => " 68_delay", delay_value => 1)  port map(req => inputPort_4_Daemon_CP_609_elements(9), ack => inputPort_4_Daemon_CP_609_elements(68), clk => clk, reset =>reset);
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	58 
    -- CP-element group 69: 	64 
    -- CP-element group 69: 	67 
    -- CP-element group 69: 	61 
    -- CP-element group 69: 	12 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	6 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_338/do_while_stmt_339/do_while_stmt_339_loop_body/$exit
      -- 
    inputPort_4_Daemon_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "inputPort_4_Daemon_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= inputPort_4_Daemon_CP_609_elements(58) & inputPort_4_Daemon_CP_609_elements(64) & inputPort_4_Daemon_CP_609_elements(67) & inputPort_4_Daemon_CP_609_elements(61) & inputPort_4_Daemon_CP_609_elements(12);
      gj_inputPort_4_Daemon_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	5 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_338/do_while_stmt_339/loop_exit/$exit
      -- CP-element group 70: 	 branch_block_stmt_338/do_while_stmt_339/loop_exit/ack
      -- 
    ack_805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_339_branch_ack_0, ack => inputPort_4_Daemon_CP_609_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	5 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_338/do_while_stmt_339/loop_taken/$exit
      -- CP-element group 71: 	 branch_block_stmt_338/do_while_stmt_339/loop_taken/ack
      -- 
    ack_809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_339_branch_ack_1, ack => inputPort_4_Daemon_CP_609_elements(71)); -- 
    -- CP-element group 72:  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	3 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	1 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_338/do_while_stmt_339/$exit
      -- 
    inputPort_4_Daemon_CP_609_elements(72) <= inputPort_4_Daemon_CP_609_elements(3);
    inputPort_4_Daemon_do_while_stmt_339_terminator_810: loop_terminator -- 
      generic map (name => " inputPort_4_Daemon_do_while_stmt_339_terminator_810", max_iterations_in_flight =>7) 
      port map(loop_body_exit => inputPort_4_Daemon_CP_609_elements(6),loop_continue => inputPort_4_Daemon_CP_609_elements(71),loop_terminate => inputPort_4_Daemon_CP_609_elements(70),loop_back => inputPort_4_Daemon_CP_609_elements(4),loop_exit => inputPort_4_Daemon_CP_609_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_341_phi_seq_682_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_4_Daemon_CP_609_elements(21);
      inputPort_4_Daemon_CP_609_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_4_Daemon_CP_609_elements(24);
      inputPort_4_Daemon_CP_609_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_4_Daemon_CP_609_elements(26);
      inputPort_4_Daemon_CP_609_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_4_Daemon_CP_609_elements(19);
      inputPort_4_Daemon_CP_609_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_4_Daemon_CP_609_elements(30);
      inputPort_4_Daemon_CP_609_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_4_Daemon_CP_609_elements(31);
      inputPort_4_Daemon_CP_609_elements(20) <= phi_mux_reqs(1);
      phi_stmt_341_phi_seq_682 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_341_phi_seq_682") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_4_Daemon_CP_609_elements(11), 
          phi_sample_ack => inputPort_4_Daemon_CP_609_elements(17), 
          phi_update_req => inputPort_4_Daemon_CP_609_elements(13), 
          phi_update_ack => inputPort_4_Daemon_CP_609_elements(18), 
          phi_mux_ack => inputPort_4_Daemon_CP_609_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_349_phi_seq_744_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= inputPort_4_Daemon_CP_609_elements(45);
      inputPort_4_Daemon_CP_609_elements(48)<= src_sample_reqs(0);
      src_sample_acks(0)  <= inputPort_4_Daemon_CP_609_elements(48);
      inputPort_4_Daemon_CP_609_elements(49)<= src_update_reqs(0);
      src_update_acks(0)  <= inputPort_4_Daemon_CP_609_elements(50);
      inputPort_4_Daemon_CP_609_elements(46) <= phi_mux_reqs(0);
      triggers(1)  <= inputPort_4_Daemon_CP_609_elements(43);
      inputPort_4_Daemon_CP_609_elements(52)<= src_sample_reqs(1);
      src_sample_acks(1)  <= inputPort_4_Daemon_CP_609_elements(54);
      inputPort_4_Daemon_CP_609_elements(53)<= src_update_reqs(1);
      src_update_acks(1)  <= inputPort_4_Daemon_CP_609_elements(55);
      inputPort_4_Daemon_CP_609_elements(44) <= phi_mux_reqs(1);
      phi_stmt_349_phi_seq_744 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_349_phi_seq_744") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => inputPort_4_Daemon_CP_609_elements(39), 
          phi_sample_ack => inputPort_4_Daemon_CP_609_elements(40), 
          phi_update_req => inputPort_4_Daemon_CP_609_elements(41), 
          phi_update_ack => inputPort_4_Daemon_CP_609_elements(42), 
          phi_mux_ack => inputPort_4_Daemon_CP_609_elements(47), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_634_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= inputPort_4_Daemon_CP_609_elements(7);
        preds(1)  <= inputPort_4_Daemon_CP_609_elements(8);
        entry_tmerge_634 : transition_merge -- 
          generic map(name => " entry_tmerge_634")
          port map (preds => preds, symbol_out => inputPort_4_Daemon_CP_609_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal RPIPE_in_data_4_348_wire : std_logic_vector(31 downto 0);
    signal R_ONE_1_384_wire_constant : std_logic_vector(0 downto 0);
    signal SUB_u16_u16_371_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_374_wire : std_logic_vector(15 downto 0);
    signal count_down_341 : std_logic_vector(15 downto 0);
    signal data_to_outport_387 : std_logic_vector(32 downto 0);
    signal dest_id_362 : std_logic_vector(7 downto 0);
    signal input_word_346 : std_logic_vector(31 downto 0);
    signal konst_351_wire_constant : std_logic_vector(7 downto 0);
    signal konst_356_wire_constant : std_logic_vector(15 downto 0);
    signal konst_370_wire_constant : std_logic_vector(15 downto 0);
    signal konst_373_wire_constant : std_logic_vector(15 downto 0);
    signal konst_390_wire_constant : std_logic_vector(7 downto 0);
    signal konst_399_wire_constant : std_logic_vector(7 downto 0);
    signal konst_408_wire_constant : std_logic_vector(7 downto 0);
    signal konst_417_wire_constant : std_logic_vector(7 downto 0);
    signal konst_425_wire_constant : std_logic_vector(0 downto 0);
    signal last_dest_id_349 : std_logic_vector(7 downto 0);
    signal new_packet_358 : std_logic_vector(0 downto 0);
    signal next_count_down_376 : std_logic_vector(15 downto 0);
    signal next_count_down_376_345_buffered : std_logic_vector(15 downto 0);
    signal next_last_dest_id_382 : std_logic_vector(7 downto 0);
    signal next_last_dest_id_382_352_buffered : std_logic_vector(7 downto 0);
    signal pkt_length_366 : std_logic_vector(15 downto 0);
    signal send_to_1_392 : std_logic_vector(0 downto 0);
    signal send_to_2_401 : std_logic_vector(0 downto 0);
    signal send_to_3_410 : std_logic_vector(0 downto 0);
    signal send_to_4_419 : std_logic_vector(0 downto 0);
    signal type_cast_344_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    R_ONE_1_384_wire_constant <= "1";
    konst_351_wire_constant <= "00000000";
    konst_356_wire_constant <= "0000000000000000";
    konst_370_wire_constant <= "0000000000000001";
    konst_373_wire_constant <= "0000000000000001";
    konst_390_wire_constant <= "00000001";
    konst_399_wire_constant <= "00000010";
    konst_408_wire_constant <= "00000011";
    konst_417_wire_constant <= "00000100";
    konst_425_wire_constant <= "1";
    type_cast_344_wire_constant <= "0000000000000000";
    phi_stmt_341: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_344_wire_constant & next_count_down_376_345_buffered;
      req <= phi_stmt_341_req_0 & phi_stmt_341_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_341",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_341_ack_0,
          idata => idata,
          odata => count_down_341,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_341
    phi_stmt_349: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_351_wire_constant & next_last_dest_id_382_352_buffered;
      req <= phi_stmt_349_req_0 & phi_stmt_349_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_349",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_349_ack_0,
          idata => idata,
          odata => last_dest_id_349,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_349
    -- flow-through select operator MUX_375_inst
    next_count_down_376 <= SUB_u16_u16_371_wire when (new_packet_358(0) /=  '0') else SUB_u16_u16_374_wire;
    -- flow-through select operator MUX_381_inst
    next_last_dest_id_382 <= dest_id_362 when (new_packet_358(0) /=  '0') else last_dest_id_349;
    -- flow-through slice operator slice_361_inst
    dest_id_362 <= input_word_346(31 downto 24);
    -- flow-through slice operator slice_365_inst
    pkt_length_366 <= input_word_346(23 downto 8);
    next_count_down_376_345_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_count_down_376_345_buf_req_0;
      next_count_down_376_345_buf_ack_0<= wack(0);
      rreq(0) <= next_count_down_376_345_buf_req_1;
      next_count_down_376_345_buf_ack_1<= rack(0);
      next_count_down_376_345_buf : InterlockBuffer generic map ( -- 
        name => "next_count_down_376_345_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_count_down_376,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_count_down_376_345_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_last_dest_id_382_352_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_last_dest_id_382_352_buf_req_0;
      next_last_dest_id_382_352_buf_ack_0<= wack(0);
      rreq(0) <= next_last_dest_id_382_352_buf_req_1;
      next_last_dest_id_382_352_buf_ack_1<= rack(0);
      next_last_dest_id_382_352_buf : InterlockBuffer generic map ( -- 
        name => "next_last_dest_id_382_352_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_last_dest_id_382,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_last_dest_id_382_352_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_346
    process(RPIPE_in_data_4_348_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := RPIPE_in_data_4_348_wire(31 downto 0);
      input_word_346 <= tmp_var; -- 
    end process;
    do_while_stmt_339_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_425_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_339_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_339_branch_req_0,
          ack0 => do_while_stmt_339_branch_ack_0,
          ack1 => do_while_stmt_339_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator CONCAT_u1_u33_386_inst
    process(R_ONE_1_384_wire_constant, input_word_346) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(R_ONE_1_384_wire_constant, input_word_346, tmp_var);
      data_to_outport_387 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_357_inst
    process(count_down_341) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(count_down_341, konst_356_wire_constant, tmp_var);
      new_packet_358 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_391_inst
    process(next_last_dest_id_382) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_382, konst_390_wire_constant, tmp_var);
      send_to_1_392 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_400_inst
    process(next_last_dest_id_382) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_382, konst_399_wire_constant, tmp_var);
      send_to_2_401 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_409_inst
    process(next_last_dest_id_382) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_382, konst_408_wire_constant, tmp_var);
      send_to_3_410 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_418_inst
    process(next_last_dest_id_382) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_last_dest_id_382, konst_417_wire_constant, tmp_var);
      send_to_4_419 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_371_inst
    process(pkt_length_366) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(pkt_length_366, konst_370_wire_constant, tmp_var);
      SUB_u16_u16_371_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_374_inst
    process(count_down_341) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(count_down_341, konst_373_wire_constant, tmp_var);
      SUB_u16_u16_374_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_in_data_4_348_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_in_data_4_348_inst_req_0;
      RPIPE_in_data_4_348_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_in_data_4_348_inst_req_1;
      RPIPE_in_data_4_348_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_in_data_4_348_wire <= data_out(31 downto 0);
      in_data_4_read_0_gI: SplitGuardInterface generic map(name => "in_data_4_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      in_data_4_read_0: InputPortRevised -- 
        generic map ( name => "in_data_4_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => in_data_4_pipe_read_req(0),
          oack => in_data_4_pipe_read_ack(0),
          odata => in_data_4_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_noblock_obuf_4_1_394_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_4_1_394_inst_req_0;
      WPIPE_noblock_obuf_4_1_394_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_4_1_394_inst_req_1;
      WPIPE_noblock_obuf_4_1_394_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_1_392(0);
      data_in <= data_to_outport_387;
      noblock_obuf_4_1_write_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_1_write_0: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_4_1", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_4_1_pipe_write_req(0),
          oack => noblock_obuf_4_1_pipe_write_ack(0),
          odata => noblock_obuf_4_1_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_noblock_obuf_4_2_403_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_4_2_403_inst_req_0;
      WPIPE_noblock_obuf_4_2_403_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_4_2_403_inst_req_1;
      WPIPE_noblock_obuf_4_2_403_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_2_401(0);
      data_in <= data_to_outport_387;
      noblock_obuf_4_2_write_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_2_write_1: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_4_2", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_4_2_pipe_write_req(0),
          oack => noblock_obuf_4_2_pipe_write_ack(0),
          odata => noblock_obuf_4_2_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_noblock_obuf_4_3_412_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_4_3_412_inst_req_0;
      WPIPE_noblock_obuf_4_3_412_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_4_3_412_inst_req_1;
      WPIPE_noblock_obuf_4_3_412_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_3_410(0);
      data_in <= data_to_outport_387;
      noblock_obuf_4_3_write_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_3_write_2: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_4_3", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_4_3_pipe_write_req(0),
          oack => noblock_obuf_4_3_pipe_write_ack(0),
          odata => noblock_obuf_4_3_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_noblock_obuf_4_4_421_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_noblock_obuf_4_4_421_inst_req_0;
      WPIPE_noblock_obuf_4_4_421_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_noblock_obuf_4_4_421_inst_req_1;
      WPIPE_noblock_obuf_4_4_421_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_4_419(0);
      data_in <= data_to_outport_387;
      noblock_obuf_4_4_write_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_4_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_4_write_3: OutputPortRevised -- 
        generic map ( name => "noblock_obuf_4_4", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => noblock_obuf_4_4_pipe_write_req(0),
          oack => noblock_obuf_4_4_pipe_write_ack(0),
          odata => noblock_obuf_4_4_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end inputPort_4_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity outputPort_1_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    noblock_obuf_4_1_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_1_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_2_1_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_1_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_1_1_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_1_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_3_1_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_1_pipe_read_data : in   std_logic_vector(32 downto 0);
    out_data_1_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_1_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity outputPort_1_Daemon;
architecture outputPort_1_Daemon_arch of outputPort_1_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal outputPort_1_Daemon_CP_814_start: Boolean;
  signal outputPort_1_Daemon_CP_814_symbol: Boolean;
  -- volatile/operator module components. 
  component prioritySelect_Volatile is -- 
    port ( -- 
      down_counter : in  std_logic_vector(7 downto 0);
      active_packet : in  std_logic_vector(2 downto 0);
      pkt_priority : in  std_logic_vector(2 downto 0);
      p1_valid : in  std_logic_vector(0 downto 0);
      p2_valid : in  std_logic_vector(0 downto 0);
      p3_valid : in  std_logic_vector(0 downto 0);
      p4_valid : in  std_logic_vector(0 downto 0);
      next_active_packet : out  std_logic_vector(2 downto 0);
      next_pkt_priority : out  std_logic_vector(2 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal do_while_stmt_655_branch_ack_1 : boolean;
  signal WPIPE_out_data_1_868_inst_ack_1 : boolean;
  signal WPIPE_out_data_1_868_inst_req_1 : boolean;
  signal WPIPE_out_data_1_868_inst_ack_0 : boolean;
  signal WPIPE_out_data_1_868_inst_req_0 : boolean;
  signal do_while_stmt_655_branch_req_0 : boolean;
  signal do_while_stmt_655_branch_ack_0 : boolean;
  signal phi_stmt_657_req_1 : boolean;
  signal phi_stmt_657_req_0 : boolean;
  signal phi_stmt_657_ack_0 : boolean;
  signal next_down_counter_772_660_buf_req_0 : boolean;
  signal next_down_counter_772_660_buf_ack_0 : boolean;
  signal next_down_counter_772_660_buf_req_1 : boolean;
  signal next_down_counter_772_660_buf_ack_1 : boolean;
  signal phi_stmt_661_req_1 : boolean;
  signal phi_stmt_661_req_0 : boolean;
  signal phi_stmt_661_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_1_665_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_1_1_665_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_1_665_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_1_1_665_inst_ack_1 : boolean;
  signal phi_stmt_666_req_1 : boolean;
  signal phi_stmt_666_req_0 : boolean;
  signal phi_stmt_666_ack_0 : boolean;
  signal RPIPE_noblock_obuf_2_1_670_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_2_1_670_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_2_1_670_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_2_1_670_inst_ack_1 : boolean;
  signal phi_stmt_671_req_1 : boolean;
  signal phi_stmt_671_req_0 : boolean;
  signal phi_stmt_671_ack_0 : boolean;
  signal RPIPE_noblock_obuf_3_1_675_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_3_1_675_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_3_1_675_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_3_1_675_inst_ack_1 : boolean;
  signal phi_stmt_676_req_1 : boolean;
  signal phi_stmt_676_req_0 : boolean;
  signal phi_stmt_676_ack_0 : boolean;
  signal RPIPE_noblock_obuf_4_1_680_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_4_1_680_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_4_1_680_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_4_1_680_inst_ack_1 : boolean;
  signal phi_stmt_681_req_1 : boolean;
  signal phi_stmt_681_req_0 : boolean;
  signal phi_stmt_681_ack_0 : boolean;
  signal next_active_packet_748_684_buf_req_0 : boolean;
  signal next_active_packet_748_684_buf_ack_0 : boolean;
  signal next_active_packet_748_684_buf_req_1 : boolean;
  signal next_active_packet_748_684_buf_ack_1 : boolean;
  signal phi_stmt_685_req_1 : boolean;
  signal phi_stmt_685_req_0 : boolean;
  signal phi_stmt_685_ack_0 : boolean;
  signal next_pkt_priority_748_688_buf_req_0 : boolean;
  signal next_pkt_priority_748_688_buf_ack_0 : boolean;
  signal next_pkt_priority_748_688_buf_req_1 : boolean;
  signal next_pkt_priority_748_688_buf_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "outputPort_1_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  outputPort_1_Daemon_CP_814_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "outputPort_1_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_1_Daemon_CP_814_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= outputPort_1_Daemon_CP_814_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_1_Daemon_CP_814_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  outputPort_1_Daemon_CP_814: Block -- control-path 
    signal outputPort_1_Daemon_CP_814_elements: BooleanArray(161 downto 0);
    -- 
  begin -- 
    outputPort_1_Daemon_CP_814_elements(0) <= outputPort_1_Daemon_CP_814_start;
    outputPort_1_Daemon_CP_814_symbol <= outputPort_1_Daemon_CP_814_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_654/do_while_stmt_655__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_654/$entry
      -- CP-element group 0: 	 branch_block_stmt_654/branch_block_stmt_654__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	161 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_654/$exit
      -- CP-element group 1: 	 branch_block_stmt_654/do_while_stmt_655__exit__
      -- CP-element group 1: 	 branch_block_stmt_654/branch_block_stmt_654__exit__
      -- CP-element group 1: 	 $exit
      -- 
    outputPort_1_Daemon_CP_814_elements(1) <= outputPort_1_Daemon_CP_814_elements(161);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_654/do_while_stmt_655/$entry
      -- CP-element group 2: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655__entry__
      -- 
    outputPort_1_Daemon_CP_814_elements(2) <= outputPort_1_Daemon_CP_814_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	161 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655__exit__
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_654/do_while_stmt_655/loop_back
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	160 
    -- CP-element group 5: 	159 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_654/do_while_stmt_655/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_654/do_while_stmt_655/condition_done
      -- CP-element group 5: 	 branch_block_stmt_654/do_while_stmt_655/loop_taken/$entry
      -- 
    outputPort_1_Daemon_CP_814_elements(5) <= outputPort_1_Daemon_CP_814_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	158 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_654/do_while_stmt_655/loop_body_done
      -- 
    outputPort_1_Daemon_CP_814_elements(6) <= outputPort_1_Daemon_CP_814_elements(158);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	141 
    -- CP-element group 7: 	102 
    -- CP-element group 7: 	122 
    -- CP-element group 7: 	21 
    -- CP-element group 7: 	40 
    -- CP-element group 7: 	61 
    -- CP-element group 7: 	82 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/back_edge_to_loop_body
      -- 
    outputPort_1_Daemon_CP_814_elements(7) <= outputPort_1_Daemon_CP_814_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	104 
    -- CP-element group 8: 	124 
    -- CP-element group 8: 	143 
    -- CP-element group 8: 	23 
    -- CP-element group 8: 	42 
    -- CP-element group 8: 	63 
    -- CP-element group 8: 	84 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/first_time_through_loop_body
      -- 
    outputPort_1_Daemon_CP_814_elements(8) <= outputPort_1_Daemon_CP_814_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	135 
    -- CP-element group 9: 	117 
    -- CP-element group 9: 	98 
    -- CP-element group 9: 	118 
    -- CP-element group 9: 	157 
    -- CP-element group 9: 	136 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	34 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	55 
    -- CP-element group 9: 	56 
    -- CP-element group 9: 	76 
    -- CP-element group 9: 	77 
    -- CP-element group 9: 	97 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/loop_body_start
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	157 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/condition_evaluated
      -- 
    condition_evaluated_838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(10), ack => do_while_stmt_655_branch_req_0); -- 
    outputPort_1_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(157) & outputPort_1_Daemon_CP_814_elements(14);
      gj_outputPort_1_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	135 
    -- CP-element group 11: 	117 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	55 
    -- CP-element group 11: 	76 
    -- CP-element group 11: 	97 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	137 
    -- CP-element group 11: 	99 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	57 
    -- CP-element group 11: 	78 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_681_sample_start__ps
      -- 
    outputPort_1_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(135) & outputPort_1_Daemon_CP_814_elements(117) & outputPort_1_Daemon_CP_814_elements(15) & outputPort_1_Daemon_CP_814_elements(34) & outputPort_1_Daemon_CP_814_elements(55) & outputPort_1_Daemon_CP_814_elements(76) & outputPort_1_Daemon_CP_814_elements(97) & outputPort_1_Daemon_CP_814_elements(14);
      gj_outputPort_1_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	100 
    -- CP-element group 12: 	119 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	37 
    -- CP-element group 12: 	138 
    -- CP-element group 12: 	58 
    -- CP-element group 12: 	79 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	158 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	135 
    -- CP-element group 12: 	117 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	34 
    -- CP-element group 12: 	55 
    -- CP-element group 12: 	76 
    -- CP-element group 12: 	97 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_657_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_661_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_666_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_671_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_676_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_681_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_685_sample_completed_
      -- 
    outputPort_1_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(100) & outputPort_1_Daemon_CP_814_elements(119) & outputPort_1_Daemon_CP_814_elements(18) & outputPort_1_Daemon_CP_814_elements(37) & outputPort_1_Daemon_CP_814_elements(138) & outputPort_1_Daemon_CP_814_elements(58) & outputPort_1_Daemon_CP_814_elements(79);
      gj_outputPort_1_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	98 
    -- CP-element group 13: 	118 
    -- CP-element group 13: 	136 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	35 
    -- CP-element group 13: 	56 
    -- CP-element group 13: 	77 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	120 
    -- CP-element group 13: 	19 
    -- CP-element group 13: 	38 
    -- CP-element group 13: 	139 
    -- CP-element group 13: 	59 
    -- CP-element group 13: 	80 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_676_update_start__ps
      -- 
    outputPort_1_Daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(98) & outputPort_1_Daemon_CP_814_elements(118) & outputPort_1_Daemon_CP_814_elements(136) & outputPort_1_Daemon_CP_814_elements(16) & outputPort_1_Daemon_CP_814_elements(35) & outputPort_1_Daemon_CP_814_elements(56) & outputPort_1_Daemon_CP_814_elements(77);
      gj_outputPort_1_Daemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	140 
    -- CP-element group 14: 	121 
    -- CP-element group 14: 	101 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	60 
    -- CP-element group 14: 	81 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/aggregated_phi_update_ack
      -- 
    outputPort_1_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(140) & outputPort_1_Daemon_CP_814_elements(121) & outputPort_1_Daemon_CP_814_elements(101) & outputPort_1_Daemon_CP_814_elements(20) & outputPort_1_Daemon_CP_814_elements(39) & outputPort_1_Daemon_CP_814_elements(60) & outputPort_1_Daemon_CP_814_elements(81);
      gj_outputPort_1_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_657_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	155 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_657_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(155);
      gj_outputPort_1_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_657_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(17) <= outputPort_1_Daemon_CP_814_elements(11);
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_657_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_657_update_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(19) <= outputPort_1_Daemon_CP_814_elements(13);
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	154 
    -- CP-element group 20: 	14 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_657_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_657_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_657_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(21) <= outputPort_1_Daemon_CP_814_elements(7);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_657_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_657_loopback_sample_req_ps
      -- 
    phi_stmt_657_loopback_sample_req_853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_657_loopback_sample_req_853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(22), ack => phi_stmt_657_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_657_entry_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(23) <= outputPort_1_Daemon_CP_814_elements(8);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_657_entry_sample_req
      -- CP-element group 24: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_657_entry_sample_req_ps
      -- 
    phi_stmt_657_entry_sample_req_856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_657_entry_sample_req_856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(24), ack => phi_stmt_657_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_657_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_657_phi_mux_ack_ps
      -- 
    phi_stmt_657_phi_mux_ack_859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_657_ack_0, ack => outputPort_1_Daemon_CP_814_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_8_659_sample_start__ps
      -- CP-element group 26: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_8_659_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_8_659_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_8_659_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_8_659_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_8_659_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_8_659_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(28) <= outputPort_1_Daemon_CP_814_elements(29);
    -- CP-element group 29:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	28 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_8_659_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(29) is a control-delay.
    cp_element_29_delay: control_delay_element  generic map(name => " 29_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_814_elements(27), ack => outputPort_1_Daemon_CP_814_elements(29), clk => clk, reset =>reset);
    -- CP-element group 30:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_down_counter_660_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_down_counter_660_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_down_counter_660_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_down_counter_660_Sample/req
      -- 
    req_880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(30), ack => next_down_counter_772_660_buf_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_down_counter_660_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_down_counter_660_update_start_
      -- CP-element group 31: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_down_counter_660_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_down_counter_660_Update/req
      -- 
    req_885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(31), ack => next_down_counter_772_660_buf_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_down_counter_660_sample_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_down_counter_660_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_down_counter_660_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_down_counter_660_Sample/ack
      -- 
    ack_881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_772_660_buf_ack_0, ack => outputPort_1_Daemon_CP_814_elements(32)); -- 
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_down_counter_660_update_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_down_counter_660_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_down_counter_660_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_down_counter_660_Update/ack
      -- 
    ack_886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_772_660_buf_ack_1, ack => outputPort_1_Daemon_CP_814_elements(33)); -- 
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	9 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	12 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	11 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_661_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	155 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	13 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_661_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(155);
      gj_outputPort_1_Daemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	11 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_661_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(36) <= outputPort_1_Daemon_CP_814_elements(11);
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	12 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_661_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_661_update_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(38) <= outputPort_1_Daemon_CP_814_elements(13);
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	154 
    -- CP-element group 39: 	14 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_661_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_661_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	7 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_661_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(40) <= outputPort_1_Daemon_CP_814_elements(7);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_661_loopback_sample_req
      -- CP-element group 41: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_661_loopback_sample_req_ps
      -- 
    phi_stmt_661_loopback_sample_req_897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_661_loopback_sample_req_897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(41), ack => phi_stmt_661_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	8 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_661_entry_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(42) <= outputPort_1_Daemon_CP_814_elements(8);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_661_entry_sample_req
      -- CP-element group 43: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_661_entry_sample_req_ps
      -- 
    phi_stmt_661_entry_sample_req_900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_661_entry_sample_req_900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(43), ack => phi_stmt_661_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_661_phi_mux_ack
      -- CP-element group 44: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_661_phi_mux_ack_ps
      -- 
    phi_stmt_661_phi_mux_ack_903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_661_ack_0, ack => outputPort_1_Daemon_CP_814_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_663_sample_start__ps
      -- CP-element group 45: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_663_sample_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_663_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_663_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_663_update_start__ps
      -- CP-element group 46: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_663_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_663_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(47) <= outputPort_1_Daemon_CP_814_elements(48);
    -- CP-element group 48:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	47 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_663_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(48) is a control-delay.
    cp_element_48_delay: control_delay_element  generic map(name => " 48_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_814_elements(46), ack => outputPort_1_Daemon_CP_814_elements(48), clk => clk, reset =>reset);
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_1_1_665_sample_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_1_1_665_update_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	54 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_1_1_665_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_1_1_665_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_1_1_665_Sample/rr
      -- 
    rr_924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(51), ack => RPIPE_noblock_obuf_1_1_665_inst_req_0); -- 
    outputPort_1_Daemon_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(49) & outputPort_1_Daemon_CP_814_elements(54);
      gj_outputPort_1_Daemon_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: 	53 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_1_1_665_update_start_
      -- CP-element group 52: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_1_1_665_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_1_1_665_Update/cr
      -- 
    cr_929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(52), ack => RPIPE_noblock_obuf_1_1_665_inst_req_1); -- 
    outputPort_1_Daemon_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(50) & outputPort_1_Daemon_CP_814_elements(53);
      gj_outputPort_1_Daemon_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	52 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_1_1_665_sample_completed__ps
      -- CP-element group 53: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_1_1_665_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_1_1_665_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_1_1_665_Sample/ra
      -- 
    ra_925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_1_665_inst_ack_0, ack => outputPort_1_Daemon_CP_814_elements(53)); -- 
    -- CP-element group 54:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	51 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_1_1_665_update_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_1_1_665_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_1_1_665_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_1_1_665_Update/ca
      -- 
    ca_930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_1_665_inst_ack_1, ack => outputPort_1_Daemon_CP_814_elements(54)); -- 
    -- CP-element group 55:  join  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	9 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	12 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	11 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_666_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	9 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	155 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	13 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_666_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(155);
      gj_outputPort_1_Daemon_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	11 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_666_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(57) <= outputPort_1_Daemon_CP_814_elements(11);
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	12 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_666_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	13 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_666_update_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(59) <= outputPort_1_Daemon_CP_814_elements(13);
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	154 
    -- CP-element group 60: 	14 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_666_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_666_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	7 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_666_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(61) <= outputPort_1_Daemon_CP_814_elements(7);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_666_loopback_sample_req
      -- CP-element group 62: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_666_loopback_sample_req_ps
      -- 
    phi_stmt_666_loopback_sample_req_941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_666_loopback_sample_req_941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(62), ack => phi_stmt_666_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	8 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_666_entry_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(63) <= outputPort_1_Daemon_CP_814_elements(8);
    -- CP-element group 64:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_666_entry_sample_req
      -- CP-element group 64: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_666_entry_sample_req_ps
      -- 
    phi_stmt_666_entry_sample_req_944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_666_entry_sample_req_944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(64), ack => phi_stmt_666_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_666_phi_mux_ack
      -- CP-element group 65: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_666_phi_mux_ack_ps
      -- 
    phi_stmt_666_phi_mux_ack_947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_666_ack_0, ack => outputPort_1_Daemon_CP_814_elements(65)); -- 
    -- CP-element group 66:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_668_sample_start__ps
      -- CP-element group 66: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_668_sample_completed__ps
      -- CP-element group 66: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_668_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_668_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_668_update_start__ps
      -- CP-element group 67: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_668_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_668_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(68) <= outputPort_1_Daemon_CP_814_elements(69);
    -- CP-element group 69:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	68 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_668_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(69) is a control-delay.
    cp_element_69_delay: control_delay_element  generic map(name => " 69_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_814_elements(67), ack => outputPort_1_Daemon_CP_814_elements(69), clk => clk, reset =>reset);
    -- CP-element group 70:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_2_1_670_sample_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(70) is bound as output of CP function.
    -- CP-element group 71:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_2_1_670_update_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: marked-predecessors 
    -- CP-element group 72: 	75 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_2_1_670_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_2_1_670_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_2_1_670_Sample/rr
      -- 
    rr_968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(72), ack => RPIPE_noblock_obuf_2_1_670_inst_req_0); -- 
    outputPort_1_Daemon_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(70) & outputPort_1_Daemon_CP_814_elements(75);
      gj_outputPort_1_Daemon_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: 	74 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_2_1_670_update_start_
      -- CP-element group 73: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_2_1_670_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_2_1_670_Update/cr
      -- 
    cr_973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(73), ack => RPIPE_noblock_obuf_2_1_670_inst_req_1); -- 
    outputPort_1_Daemon_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(71) & outputPort_1_Daemon_CP_814_elements(74);
      gj_outputPort_1_Daemon_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	73 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_2_1_670_sample_completed__ps
      -- CP-element group 74: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_2_1_670_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_2_1_670_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_2_1_670_Sample/ra
      -- 
    ra_969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_1_670_inst_ack_0, ack => outputPort_1_Daemon_CP_814_elements(74)); -- 
    -- CP-element group 75:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	72 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_2_1_670_update_completed__ps
      -- CP-element group 75: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_2_1_670_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_2_1_670_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_2_1_670_Update/ca
      -- 
    ca_974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_1_670_inst_ack_1, ack => outputPort_1_Daemon_CP_814_elements(75)); -- 
    -- CP-element group 76:  join  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	9 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	12 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	11 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_671_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	9 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	155 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	13 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_671_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(155);
      gj_outputPort_1_Daemon_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	11 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_671_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(78) <= outputPort_1_Daemon_CP_814_elements(11);
    -- CP-element group 79:  join  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	12 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_671_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	13 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_671_update_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(80) <= outputPort_1_Daemon_CP_814_elements(13);
    -- CP-element group 81:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	154 
    -- CP-element group 81: 	14 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_671_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_671_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	7 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_671_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(82) <= outputPort_1_Daemon_CP_814_elements(7);
    -- CP-element group 83:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_671_loopback_sample_req
      -- CP-element group 83: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_671_loopback_sample_req_ps
      -- 
    phi_stmt_671_loopback_sample_req_985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_671_loopback_sample_req_985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(83), ack => phi_stmt_671_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(83) is bound as output of CP function.
    -- CP-element group 84:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	8 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_671_entry_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(84) <= outputPort_1_Daemon_CP_814_elements(8);
    -- CP-element group 85:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_671_entry_sample_req
      -- CP-element group 85: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_671_entry_sample_req_ps
      -- 
    phi_stmt_671_entry_sample_req_988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_671_entry_sample_req_988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(85), ack => phi_stmt_671_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_671_phi_mux_ack_ps
      -- CP-element group 86: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_671_phi_mux_ack
      -- 
    phi_stmt_671_phi_mux_ack_991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_671_ack_0, ack => outputPort_1_Daemon_CP_814_elements(86)); -- 
    -- CP-element group 87:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_673_sample_start__ps
      -- CP-element group 87: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_673_sample_completed__ps
      -- CP-element group 87: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_673_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_673_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_673_update_start__ps
      -- CP-element group 88: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_673_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	90 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_673_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(89) <= outputPort_1_Daemon_CP_814_elements(90);
    -- CP-element group 90:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	89 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_673_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(90) is a control-delay.
    cp_element_90_delay: control_delay_element  generic map(name => " 90_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_814_elements(88), ack => outputPort_1_Daemon_CP_814_elements(90), clk => clk, reset =>reset);
    -- CP-element group 91:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_3_1_675_sample_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(91) is bound as output of CP function.
    -- CP-element group 92:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_3_1_675_update_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(92) is bound as output of CP function.
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	96 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_3_1_675_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_3_1_675_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_3_1_675_Sample/rr
      -- 
    rr_1012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(93), ack => RPIPE_noblock_obuf_3_1_675_inst_req_0); -- 
    outputPort_1_Daemon_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(91) & outputPort_1_Daemon_CP_814_elements(96);
      gj_outputPort_1_Daemon_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	95 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_3_1_675_update_start_
      -- CP-element group 94: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_3_1_675_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_3_1_675_Update/cr
      -- 
    cr_1017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(94), ack => RPIPE_noblock_obuf_3_1_675_inst_req_1); -- 
    outputPort_1_Daemon_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(92) & outputPort_1_Daemon_CP_814_elements(95);
      gj_outputPort_1_Daemon_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	94 
    -- CP-element group 95:  members (4) 
      -- CP-element group 95: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_3_1_675_sample_completed__ps
      -- CP-element group 95: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_3_1_675_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_3_1_675_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_3_1_675_Sample/ra
      -- 
    ra_1013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_1_675_inst_ack_0, ack => outputPort_1_Daemon_CP_814_elements(95)); -- 
    -- CP-element group 96:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	93 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_3_1_675_update_completed__ps
      -- CP-element group 96: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_3_1_675_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_3_1_675_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_3_1_675_Update/ca
      -- 
    ca_1018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_1_675_inst_ack_1, ack => outputPort_1_Daemon_CP_814_elements(96)); -- 
    -- CP-element group 97:  join  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	9 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	12 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	11 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_676_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	9 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	155 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	13 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_676_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_1_Daemon_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(155);
      gj_outputPort_1_Daemon_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	11 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_676_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(99) <= outputPort_1_Daemon_CP_814_elements(11);
    -- CP-element group 100:  join  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	12 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_676_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(100) is bound as output of CP function.
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	154 
    -- CP-element group 101: 	14 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_676_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_676_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(101) is bound as output of CP function.
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	7 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_676_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(102) <= outputPort_1_Daemon_CP_814_elements(7);
    -- CP-element group 103:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_676_loopback_sample_req
      -- CP-element group 103: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_676_loopback_sample_req_ps
      -- 
    phi_stmt_676_loopback_sample_req_1029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_676_loopback_sample_req_1029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(103), ack => phi_stmt_676_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(103) is bound as output of CP function.
    -- CP-element group 104:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	8 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_676_entry_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(104) <= outputPort_1_Daemon_CP_814_elements(8);
    -- CP-element group 105:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_676_entry_sample_req
      -- CP-element group 105: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_676_entry_sample_req_ps
      -- 
    phi_stmt_676_entry_sample_req_1032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_676_entry_sample_req_1032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(105), ack => phi_stmt_676_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(105) is bound as output of CP function.
    -- CP-element group 106:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_676_phi_mux_ack
      -- CP-element group 106: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_676_phi_mux_ack_ps
      -- 
    phi_stmt_676_phi_mux_ack_1035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_676_ack_0, ack => outputPort_1_Daemon_CP_814_elements(106)); -- 
    -- CP-element group 107:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (4) 
      -- CP-element group 107: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_678_sample_start__ps
      -- CP-element group 107: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_678_sample_completed__ps
      -- CP-element group 107: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_678_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_678_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(107) is bound as output of CP function.
    -- CP-element group 108:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_678_update_start__ps
      -- CP-element group 108: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_678_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(108) is bound as output of CP function.
    -- CP-element group 109:  join  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	110 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_678_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(109) <= outputPort_1_Daemon_CP_814_elements(110);
    -- CP-element group 110:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	109 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_33_678_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(110) is a control-delay.
    cp_element_110_delay: control_delay_element  generic map(name => " 110_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_814_elements(108), ack => outputPort_1_Daemon_CP_814_elements(110), clk => clk, reset =>reset);
    -- CP-element group 111:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_4_1_680_sample_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(111) is bound as output of CP function.
    -- CP-element group 112:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_4_1_680_update_start__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(112) is bound as output of CP function.
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	116 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_4_1_680_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_4_1_680_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_4_1_680_Sample/rr
      -- 
    rr_1056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(113), ack => RPIPE_noblock_obuf_4_1_680_inst_req_0); -- 
    outputPort_1_Daemon_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(111) & outputPort_1_Daemon_CP_814_elements(116);
      gj_outputPort_1_Daemon_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	115 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_4_1_680_update_start_
      -- CP-element group 114: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_4_1_680_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_4_1_680_Update/cr
      -- 
    cr_1061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(114), ack => RPIPE_noblock_obuf_4_1_680_inst_req_1); -- 
    outputPort_1_Daemon_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(115) & outputPort_1_Daemon_CP_814_elements(112);
      gj_outputPort_1_Daemon_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	114 
    -- CP-element group 115:  members (4) 
      -- CP-element group 115: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_4_1_680_sample_completed__ps
      -- CP-element group 115: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_4_1_680_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_4_1_680_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_4_1_680_Sample/ra
      -- 
    ra_1057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_1_680_inst_ack_0, ack => outputPort_1_Daemon_CP_814_elements(115)); -- 
    -- CP-element group 116:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: marked-successors 
    -- CP-element group 116: 	113 
    -- CP-element group 116:  members (4) 
      -- CP-element group 116: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_4_1_680_update_completed__ps
      -- CP-element group 116: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_4_1_680_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_4_1_680_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/RPIPE_noblock_obuf_4_1_680_Update/ca
      -- 
    ca_1062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_1_680_inst_ack_1, ack => outputPort_1_Daemon_CP_814_elements(116)); -- 
    -- CP-element group 117:  join  transition  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	9 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	12 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	11 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_681_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	9 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	155 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	13 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_681_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(155);
      gj_outputPort_1_Daemon_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  join  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	12 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_681_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(119) is bound as output of CP function.
    -- CP-element group 120:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	13 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_681_update_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(120) <= outputPort_1_Daemon_CP_814_elements(13);
    -- CP-element group 121:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	154 
    -- CP-element group 121: 	14 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_681_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_681_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(121) is bound as output of CP function.
    -- CP-element group 122:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	7 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_681_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(122) <= outputPort_1_Daemon_CP_814_elements(7);
    -- CP-element group 123:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_681_loopback_sample_req
      -- CP-element group 123: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_681_loopback_sample_req_ps
      -- 
    phi_stmt_681_loopback_sample_req_1073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_681_loopback_sample_req_1073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(123), ack => phi_stmt_681_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(123) is bound as output of CP function.
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	8 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_681_entry_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(124) <= outputPort_1_Daemon_CP_814_elements(8);
    -- CP-element group 125:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_681_entry_sample_req
      -- CP-element group 125: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_681_entry_sample_req_ps
      -- 
    phi_stmt_681_entry_sample_req_1076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_681_entry_sample_req_1076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(125), ack => phi_stmt_681_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(125) is bound as output of CP function.
    -- CP-element group 126:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_681_phi_mux_ack
      -- CP-element group 126: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_681_phi_mux_ack_ps
      -- 
    phi_stmt_681_phi_mux_ack_1079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_681_ack_0, ack => outputPort_1_Daemon_CP_814_elements(126)); -- 
    -- CP-element group 127:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (4) 
      -- CP-element group 127: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_3_683_sample_start__ps
      -- CP-element group 127: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_3_683_sample_completed__ps
      -- CP-element group 127: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_3_683_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_3_683_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(127) is bound as output of CP function.
    -- CP-element group 128:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_3_683_update_start__ps
      -- CP-element group 128: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_3_683_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(128) is bound as output of CP function.
    -- CP-element group 129:  join  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	130 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_3_683_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(129) <= outputPort_1_Daemon_CP_814_elements(130);
    -- CP-element group 130:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	129 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_3_683_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(130) is a control-delay.
    cp_element_130_delay: control_delay_element  generic map(name => " 130_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_814_elements(128), ack => outputPort_1_Daemon_CP_814_elements(130), clk => clk, reset =>reset);
    -- CP-element group 131:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (4) 
      -- CP-element group 131: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_active_packet_684_sample_start__ps
      -- CP-element group 131: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_active_packet_684_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_active_packet_684_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_active_packet_684_Sample/req
      -- 
    req_1100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(131), ack => next_active_packet_748_684_buf_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(131) is bound as output of CP function.
    -- CP-element group 132:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (4) 
      -- CP-element group 132: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_active_packet_684_update_start__ps
      -- CP-element group 132: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_active_packet_684_update_start_
      -- CP-element group 132: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_active_packet_684_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_active_packet_684_Update/req
      -- 
    req_1105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(132), ack => next_active_packet_748_684_buf_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(132) is bound as output of CP function.
    -- CP-element group 133:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_active_packet_684_sample_completed__ps
      -- CP-element group 133: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_active_packet_684_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_active_packet_684_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_active_packet_684_Sample/ack
      -- 
    ack_1101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_748_684_buf_ack_0, ack => outputPort_1_Daemon_CP_814_elements(133)); -- 
    -- CP-element group 134:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_active_packet_684_update_completed__ps
      -- CP-element group 134: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_active_packet_684_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_active_packet_684_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_active_packet_684_Update/ack
      -- 
    ack_1106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_748_684_buf_ack_1, ack => outputPort_1_Daemon_CP_814_elements(134)); -- 
    -- CP-element group 135:  join  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	9 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	12 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	11 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_685_sample_start_
      -- 
    outputPort_1_Daemon_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	9 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	155 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	13 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_685_update_start_
      -- 
    outputPort_1_Daemon_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(9) & outputPort_1_Daemon_CP_814_elements(155);
      gj_outputPort_1_Daemon_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	11 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_685_sample_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(137) <= outputPort_1_Daemon_CP_814_elements(11);
    -- CP-element group 138:  join  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	12 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_685_sample_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(138) is bound as output of CP function.
    -- CP-element group 139:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	13 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_685_update_start__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(139) <= outputPort_1_Daemon_CP_814_elements(13);
    -- CP-element group 140:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	154 
    -- CP-element group 140: 	14 
    -- CP-element group 140:  members (2) 
      -- CP-element group 140: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_685_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_685_update_completed__ps
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(140) is bound as output of CP function.
    -- CP-element group 141:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	7 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_685_loopback_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(141) <= outputPort_1_Daemon_CP_814_elements(7);
    -- CP-element group 142:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_685_loopback_sample_req
      -- CP-element group 142: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_685_loopback_sample_req_ps
      -- 
    phi_stmt_685_loopback_sample_req_1117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_685_loopback_sample_req_1117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(142), ack => phi_stmt_685_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(142) is bound as output of CP function.
    -- CP-element group 143:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	8 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_685_entry_trigger
      -- 
    outputPort_1_Daemon_CP_814_elements(143) <= outputPort_1_Daemon_CP_814_elements(8);
    -- CP-element group 144:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_685_entry_sample_req
      -- CP-element group 144: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_685_entry_sample_req_ps
      -- 
    phi_stmt_685_entry_sample_req_1120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_685_entry_sample_req_1120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(144), ack => phi_stmt_685_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_685_phi_mux_ack
      -- CP-element group 145: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/phi_stmt_685_phi_mux_ack_ps
      -- 
    phi_stmt_685_phi_mux_ack_1123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_685_ack_0, ack => outputPort_1_Daemon_CP_814_elements(145)); -- 
    -- CP-element group 146:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (4) 
      -- CP-element group 146: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_3_687_sample_start__ps
      -- CP-element group 146: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_3_687_sample_completed__ps
      -- CP-element group 146: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_3_687_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_3_687_sample_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(146) is bound as output of CP function.
    -- CP-element group 147:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (2) 
      -- CP-element group 147: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_3_687_update_start__ps
      -- CP-element group 147: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_3_687_update_start_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(147) is bound as output of CP function.
    -- CP-element group 148:  join  transition  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	149 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (1) 
      -- CP-element group 148: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_3_687_update_completed__ps
      -- 
    outputPort_1_Daemon_CP_814_elements(148) <= outputPort_1_Daemon_CP_814_elements(149);
    -- CP-element group 149:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	148 
    -- CP-element group 149:  members (1) 
      -- CP-element group 149: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_ZERO_3_687_update_completed_
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(149) is a control-delay.
    cp_element_149_delay: control_delay_element  generic map(name => " 149_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_814_elements(147), ack => outputPort_1_Daemon_CP_814_elements(149), clk => clk, reset =>reset);
    -- CP-element group 150:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (4) 
      -- CP-element group 150: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_pkt_priority_688_sample_start__ps
      -- CP-element group 150: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_pkt_priority_688_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_pkt_priority_688_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_pkt_priority_688_Sample/req
      -- 
    req_1144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(150), ack => next_pkt_priority_748_688_buf_req_0); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(150) is bound as output of CP function.
    -- CP-element group 151:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (4) 
      -- CP-element group 151: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_pkt_priority_688_update_start__ps
      -- CP-element group 151: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_pkt_priority_688_update_start_
      -- CP-element group 151: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_pkt_priority_688_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_pkt_priority_688_Update/req
      -- 
    req_1149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(151), ack => next_pkt_priority_748_688_buf_req_1); -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(151) is bound as output of CP function.
    -- CP-element group 152:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (4) 
      -- CP-element group 152: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_pkt_priority_688_sample_completed__ps
      -- CP-element group 152: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_pkt_priority_688_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_pkt_priority_688_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_pkt_priority_688_Sample/ack
      -- 
    ack_1145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pkt_priority_748_688_buf_ack_0, ack => outputPort_1_Daemon_CP_814_elements(152)); -- 
    -- CP-element group 153:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (4) 
      -- CP-element group 153: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_pkt_priority_688_update_completed__ps
      -- CP-element group 153: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_pkt_priority_688_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_pkt_priority_688_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/R_next_pkt_priority_688_Update/ack
      -- 
    ack_1150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pkt_priority_748_688_buf_ack_1, ack => outputPort_1_Daemon_CP_814_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	140 
    -- CP-element group 154: 	121 
    -- CP-element group 154: 	101 
    -- CP-element group 154: 	20 
    -- CP-element group 154: 	39 
    -- CP-element group 154: 	60 
    -- CP-element group 154: 	81 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/WPIPE_out_data_1_868_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/WPIPE_out_data_1_868_Sample/req
      -- CP-element group 154: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/WPIPE_out_data_1_868_sample_start_
      -- 
    req_1159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(154), ack => WPIPE_out_data_1_868_inst_req_0); -- 
    outputPort_1_Daemon_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(140) & outputPort_1_Daemon_CP_814_elements(121) & outputPort_1_Daemon_CP_814_elements(101) & outputPort_1_Daemon_CP_814_elements(20) & outputPort_1_Daemon_CP_814_elements(39) & outputPort_1_Daemon_CP_814_elements(60) & outputPort_1_Daemon_CP_814_elements(81) & outputPort_1_Daemon_CP_814_elements(156);
      gj_outputPort_1_Daemon_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	98 
    -- CP-element group 155: 	118 
    -- CP-element group 155: 	136 
    -- CP-element group 155: 	16 
    -- CP-element group 155: 	35 
    -- CP-element group 155: 	56 
    -- CP-element group 155: 	77 
    -- CP-element group 155:  members (6) 
      -- CP-element group 155: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/WPIPE_out_data_1_868_Update/req
      -- CP-element group 155: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/WPIPE_out_data_1_868_Sample/ack
      -- CP-element group 155: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/WPIPE_out_data_1_868_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/WPIPE_out_data_1_868_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/WPIPE_out_data_1_868_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/WPIPE_out_data_1_868_update_start_
      -- 
    ack_1160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_1_868_inst_ack_0, ack => outputPort_1_Daemon_CP_814_elements(155)); -- 
    req_1164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_1_Daemon_CP_814_elements(155), ack => WPIPE_out_data_1_868_inst_req_1); -- 
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	154 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/WPIPE_out_data_1_868_Update/ack
      -- CP-element group 156: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/WPIPE_out_data_1_868_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/WPIPE_out_data_1_868_update_completed_
      -- 
    ack_1165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_1_868_inst_ack_1, ack => outputPort_1_Daemon_CP_814_elements(156)); -- 
    -- CP-element group 157:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	9 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	10 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group outputPort_1_Daemon_CP_814_elements(157) is a control-delay.
    cp_element_157_delay: control_delay_element  generic map(name => " 157_delay", delay_value => 1)  port map(req => outputPort_1_Daemon_CP_814_elements(9), ack => outputPort_1_Daemon_CP_814_elements(157), clk => clk, reset =>reset);
    -- CP-element group 158:  join  transition  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: 	12 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	6 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_654/do_while_stmt_655/do_while_stmt_655_loop_body/$exit
      -- 
    outputPort_1_Daemon_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_1_Daemon_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_1_Daemon_CP_814_elements(156) & outputPort_1_Daemon_CP_814_elements(12);
      gj_outputPort_1_Daemon_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	5 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (2) 
      -- CP-element group 159: 	 branch_block_stmt_654/do_while_stmt_655/loop_exit/$exit
      -- CP-element group 159: 	 branch_block_stmt_654/do_while_stmt_655/loop_exit/ack
      -- 
    ack_1170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_655_branch_ack_0, ack => outputPort_1_Daemon_CP_814_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	5 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (2) 
      -- CP-element group 160: 	 branch_block_stmt_654/do_while_stmt_655/loop_taken/ack
      -- CP-element group 160: 	 branch_block_stmt_654/do_while_stmt_655/loop_taken/$exit
      -- 
    ack_1174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_655_branch_ack_1, ack => outputPort_1_Daemon_CP_814_elements(160)); -- 
    -- CP-element group 161:  transition  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	3 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	1 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_654/do_while_stmt_655/$exit
      -- 
    outputPort_1_Daemon_CP_814_elements(161) <= outputPort_1_Daemon_CP_814_elements(3);
    outputPort_1_Daemon_do_while_stmt_655_terminator_1175: loop_terminator -- 
      generic map (name => " outputPort_1_Daemon_do_while_stmt_655_terminator_1175", max_iterations_in_flight =>7) 
      port map(loop_body_exit => outputPort_1_Daemon_CP_814_elements(6),loop_continue => outputPort_1_Daemon_CP_814_elements(160),loop_terminate => outputPort_1_Daemon_CP_814_elements(159),loop_back => outputPort_1_Daemon_CP_814_elements(4),loop_exit => outputPort_1_Daemon_CP_814_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_657_phi_seq_887_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_814_elements(23);
      outputPort_1_Daemon_CP_814_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_814_elements(26);
      outputPort_1_Daemon_CP_814_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_814_elements(28);
      outputPort_1_Daemon_CP_814_elements(24) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_814_elements(21);
      outputPort_1_Daemon_CP_814_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_814_elements(32);
      outputPort_1_Daemon_CP_814_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_814_elements(33);
      outputPort_1_Daemon_CP_814_elements(22) <= phi_mux_reqs(1);
      phi_stmt_657_phi_seq_887 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_657_phi_seq_887") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_814_elements(17), 
          phi_sample_ack => outputPort_1_Daemon_CP_814_elements(18), 
          phi_update_req => outputPort_1_Daemon_CP_814_elements(19), 
          phi_update_ack => outputPort_1_Daemon_CP_814_elements(20), 
          phi_mux_ack => outputPort_1_Daemon_CP_814_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_661_phi_seq_931_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_814_elements(42);
      outputPort_1_Daemon_CP_814_elements(45)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_814_elements(45);
      outputPort_1_Daemon_CP_814_elements(46)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_814_elements(47);
      outputPort_1_Daemon_CP_814_elements(43) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_814_elements(40);
      outputPort_1_Daemon_CP_814_elements(49)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_814_elements(53);
      outputPort_1_Daemon_CP_814_elements(50)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_814_elements(54);
      outputPort_1_Daemon_CP_814_elements(41) <= phi_mux_reqs(1);
      phi_stmt_661_phi_seq_931 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_661_phi_seq_931") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_814_elements(36), 
          phi_sample_ack => outputPort_1_Daemon_CP_814_elements(37), 
          phi_update_req => outputPort_1_Daemon_CP_814_elements(38), 
          phi_update_ack => outputPort_1_Daemon_CP_814_elements(39), 
          phi_mux_ack => outputPort_1_Daemon_CP_814_elements(44), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_666_phi_seq_975_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_814_elements(63);
      outputPort_1_Daemon_CP_814_elements(66)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_814_elements(66);
      outputPort_1_Daemon_CP_814_elements(67)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_814_elements(68);
      outputPort_1_Daemon_CP_814_elements(64) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_814_elements(61);
      outputPort_1_Daemon_CP_814_elements(70)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_814_elements(74);
      outputPort_1_Daemon_CP_814_elements(71)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_814_elements(75);
      outputPort_1_Daemon_CP_814_elements(62) <= phi_mux_reqs(1);
      phi_stmt_666_phi_seq_975 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_666_phi_seq_975") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_814_elements(57), 
          phi_sample_ack => outputPort_1_Daemon_CP_814_elements(58), 
          phi_update_req => outputPort_1_Daemon_CP_814_elements(59), 
          phi_update_ack => outputPort_1_Daemon_CP_814_elements(60), 
          phi_mux_ack => outputPort_1_Daemon_CP_814_elements(65), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_671_phi_seq_1019_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_814_elements(84);
      outputPort_1_Daemon_CP_814_elements(87)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_814_elements(87);
      outputPort_1_Daemon_CP_814_elements(88)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_814_elements(89);
      outputPort_1_Daemon_CP_814_elements(85) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_814_elements(82);
      outputPort_1_Daemon_CP_814_elements(91)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_814_elements(95);
      outputPort_1_Daemon_CP_814_elements(92)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_814_elements(96);
      outputPort_1_Daemon_CP_814_elements(83) <= phi_mux_reqs(1);
      phi_stmt_671_phi_seq_1019 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_671_phi_seq_1019") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_814_elements(78), 
          phi_sample_ack => outputPort_1_Daemon_CP_814_elements(79), 
          phi_update_req => outputPort_1_Daemon_CP_814_elements(80), 
          phi_update_ack => outputPort_1_Daemon_CP_814_elements(81), 
          phi_mux_ack => outputPort_1_Daemon_CP_814_elements(86), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_676_phi_seq_1063_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_814_elements(104);
      outputPort_1_Daemon_CP_814_elements(107)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_814_elements(107);
      outputPort_1_Daemon_CP_814_elements(108)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_814_elements(109);
      outputPort_1_Daemon_CP_814_elements(105) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_814_elements(102);
      outputPort_1_Daemon_CP_814_elements(111)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_814_elements(115);
      outputPort_1_Daemon_CP_814_elements(112)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_814_elements(116);
      outputPort_1_Daemon_CP_814_elements(103) <= phi_mux_reqs(1);
      phi_stmt_676_phi_seq_1063 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_676_phi_seq_1063") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_814_elements(99), 
          phi_sample_ack => outputPort_1_Daemon_CP_814_elements(100), 
          phi_update_req => outputPort_1_Daemon_CP_814_elements(13), 
          phi_update_ack => outputPort_1_Daemon_CP_814_elements(101), 
          phi_mux_ack => outputPort_1_Daemon_CP_814_elements(106), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_681_phi_seq_1107_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_814_elements(124);
      outputPort_1_Daemon_CP_814_elements(127)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_814_elements(127);
      outputPort_1_Daemon_CP_814_elements(128)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_814_elements(129);
      outputPort_1_Daemon_CP_814_elements(125) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_814_elements(122);
      outputPort_1_Daemon_CP_814_elements(131)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_814_elements(133);
      outputPort_1_Daemon_CP_814_elements(132)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_814_elements(134);
      outputPort_1_Daemon_CP_814_elements(123) <= phi_mux_reqs(1);
      phi_stmt_681_phi_seq_1107 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_681_phi_seq_1107") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_814_elements(11), 
          phi_sample_ack => outputPort_1_Daemon_CP_814_elements(119), 
          phi_update_req => outputPort_1_Daemon_CP_814_elements(120), 
          phi_update_ack => outputPort_1_Daemon_CP_814_elements(121), 
          phi_mux_ack => outputPort_1_Daemon_CP_814_elements(126), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_685_phi_seq_1151_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_1_Daemon_CP_814_elements(143);
      outputPort_1_Daemon_CP_814_elements(146)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_1_Daemon_CP_814_elements(146);
      outputPort_1_Daemon_CP_814_elements(147)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_1_Daemon_CP_814_elements(148);
      outputPort_1_Daemon_CP_814_elements(144) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_1_Daemon_CP_814_elements(141);
      outputPort_1_Daemon_CP_814_elements(150)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_1_Daemon_CP_814_elements(152);
      outputPort_1_Daemon_CP_814_elements(151)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_1_Daemon_CP_814_elements(153);
      outputPort_1_Daemon_CP_814_elements(142) <= phi_mux_reqs(1);
      phi_stmt_685_phi_seq_1151 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_685_phi_seq_1151") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_1_Daemon_CP_814_elements(137), 
          phi_sample_ack => outputPort_1_Daemon_CP_814_elements(138), 
          phi_update_req => outputPort_1_Daemon_CP_814_elements(139), 
          phi_update_ack => outputPort_1_Daemon_CP_814_elements(140), 
          phi_mux_ack => outputPort_1_Daemon_CP_814_elements(145), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_839_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= outputPort_1_Daemon_CP_814_elements(7);
        preds(1)  <= outputPort_1_Daemon_CP_814_elements(8);
        entry_tmerge_839 : transition_merge -- 
          generic map(name => " entry_tmerge_839")
          port map (preds => preds, symbol_out => outputPort_1_Daemon_CP_814_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u3_u1_713_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_719_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_726_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_732_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_778_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_786_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_794_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_802_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_808_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_815_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_823_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_830_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_841_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_847_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_854_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_860_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_759_wire : std_logic_vector(0 downto 0);
    signal MUX_716_wire : std_logic_vector(0 downto 0);
    signal MUX_722_wire : std_logic_vector(0 downto 0);
    signal MUX_729_wire : std_logic_vector(0 downto 0);
    signal MUX_735_wire : std_logic_vector(0 downto 0);
    signal MUX_770_wire : std_logic_vector(7 downto 0);
    signal MUX_812_wire : std_logic_vector(31 downto 0);
    signal MUX_819_wire : std_logic_vector(31 downto 0);
    signal MUX_827_wire : std_logic_vector(31 downto 0);
    signal MUX_834_wire : std_logic_vector(31 downto 0);
    signal MUX_844_wire : std_logic_vector(0 downto 0);
    signal MUX_850_wire : std_logic_vector(0 downto 0);
    signal MUX_857_wire : std_logic_vector(0 downto 0);
    signal MUX_863_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_775_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_783_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_791_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_799_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_723_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_736_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_752_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_755_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_756_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_851_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_864_wire : std_logic_vector(0 downto 0);
    signal OR_u32_u32_820_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_835_wire : std_logic_vector(31 downto 0);
    signal RPIPE_noblock_obuf_1_1_665_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_2_1_670_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_3_1_675_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_4_1_680_wire : std_logic_vector(32 downto 0);
    signal R_ZERO_33_663_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_668_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_673_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_678_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_3_683_wire_constant : std_logic_vector(2 downto 0);
    signal R_ZERO_3_687_wire_constant : std_logic_vector(2 downto 0);
    signal R_ZERO_8_659_wire_constant : std_logic_vector(7 downto 0);
    signal SUB_u8_u8_768_wire : std_logic_vector(7 downto 0);
    signal active_packet_681 : std_logic_vector(2 downto 0);
    signal data_to_out_837 : std_logic_vector(31 downto 0);
    signal down_counter_657 : std_logic_vector(7 downto 0);
    signal konst_692_wire_constant : std_logic_vector(32 downto 0);
    signal konst_697_wire_constant : std_logic_vector(32 downto 0);
    signal konst_702_wire_constant : std_logic_vector(32 downto 0);
    signal konst_707_wire_constant : std_logic_vector(32 downto 0);
    signal konst_712_wire_constant : std_logic_vector(2 downto 0);
    signal konst_715_wire_constant : std_logic_vector(0 downto 0);
    signal konst_718_wire_constant : std_logic_vector(2 downto 0);
    signal konst_721_wire_constant : std_logic_vector(0 downto 0);
    signal konst_725_wire_constant : std_logic_vector(2 downto 0);
    signal konst_728_wire_constant : std_logic_vector(0 downto 0);
    signal konst_731_wire_constant : std_logic_vector(2 downto 0);
    signal konst_734_wire_constant : std_logic_vector(0 downto 0);
    signal konst_758_wire_constant : std_logic_vector(7 downto 0);
    signal konst_764_wire_constant : std_logic_vector(7 downto 0);
    signal konst_767_wire_constant : std_logic_vector(7 downto 0);
    signal konst_777_wire_constant : std_logic_vector(2 downto 0);
    signal konst_785_wire_constant : std_logic_vector(2 downto 0);
    signal konst_793_wire_constant : std_logic_vector(2 downto 0);
    signal konst_801_wire_constant : std_logic_vector(2 downto 0);
    signal konst_807_wire_constant : std_logic_vector(2 downto 0);
    signal konst_811_wire_constant : std_logic_vector(31 downto 0);
    signal konst_814_wire_constant : std_logic_vector(2 downto 0);
    signal konst_818_wire_constant : std_logic_vector(31 downto 0);
    signal konst_822_wire_constant : std_logic_vector(2 downto 0);
    signal konst_826_wire_constant : std_logic_vector(31 downto 0);
    signal konst_829_wire_constant : std_logic_vector(2 downto 0);
    signal konst_833_wire_constant : std_logic_vector(31 downto 0);
    signal konst_840_wire_constant : std_logic_vector(2 downto 0);
    signal konst_843_wire_constant : std_logic_vector(0 downto 0);
    signal konst_846_wire_constant : std_logic_vector(2 downto 0);
    signal konst_849_wire_constant : std_logic_vector(0 downto 0);
    signal konst_853_wire_constant : std_logic_vector(2 downto 0);
    signal konst_856_wire_constant : std_logic_vector(0 downto 0);
    signal konst_859_wire_constant : std_logic_vector(2 downto 0);
    signal konst_862_wire_constant : std_logic_vector(0 downto 0);
    signal konst_872_wire_constant : std_logic_vector(0 downto 0);
    signal next_active_packet_748 : std_logic_vector(2 downto 0);
    signal next_active_packet_748_684_buffered : std_logic_vector(2 downto 0);
    signal next_down_counter_772 : std_logic_vector(7 downto 0);
    signal next_down_counter_772_660_buffered : std_logic_vector(7 downto 0);
    signal next_pkt_priority_748 : std_logic_vector(2 downto 0);
    signal next_pkt_priority_748_688_buffered : std_logic_vector(2 downto 0);
    signal p1_valid_694 : std_logic_vector(0 downto 0);
    signal p2_valid_699 : std_logic_vector(0 downto 0);
    signal p3_valid_704 : std_logic_vector(0 downto 0);
    signal p4_valid_709 : std_logic_vector(0 downto 0);
    signal pkt_1_e_word_661 : std_logic_vector(32 downto 0);
    signal pkt_2_e_word_666 : std_logic_vector(32 downto 0);
    signal pkt_3_e_word_671 : std_logic_vector(32 downto 0);
    signal pkt_4_e_word_676 : std_logic_vector(32 downto 0);
    signal pkt_priority_685 : std_logic_vector(2 downto 0);
    signal read_from_1_780 : std_logic_vector(0 downto 0);
    signal read_from_2_788 : std_logic_vector(0 downto 0);
    signal read_from_3_796 : std_logic_vector(0 downto 0);
    signal read_from_4_804 : std_logic_vector(0 downto 0);
    signal send_flag_866 : std_logic_vector(0 downto 0);
    signal slice_810_wire : std_logic_vector(31 downto 0);
    signal slice_817_wire : std_logic_vector(31 downto 0);
    signal slice_825_wire : std_logic_vector(31 downto 0);
    signal slice_832_wire : std_logic_vector(31 downto 0);
    signal started_new_packet_761 : std_logic_vector(0 downto 0);
    signal valid_active_pkt_word_read_738 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_ZERO_33_663_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_668_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_673_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_678_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_3_683_wire_constant <= "000";
    R_ZERO_3_687_wire_constant <= "000";
    R_ZERO_8_659_wire_constant <= "00000000";
    konst_692_wire_constant <= "000000000000000000000000000100000";
    konst_697_wire_constant <= "000000000000000000000000000100000";
    konst_702_wire_constant <= "000000000000000000000000000100000";
    konst_707_wire_constant <= "000000000000000000000000000100000";
    konst_712_wire_constant <= "001";
    konst_715_wire_constant <= "0";
    konst_718_wire_constant <= "010";
    konst_721_wire_constant <= "0";
    konst_725_wire_constant <= "011";
    konst_728_wire_constant <= "0";
    konst_731_wire_constant <= "100";
    konst_734_wire_constant <= "0";
    konst_758_wire_constant <= "00000000";
    konst_764_wire_constant <= "00111111";
    konst_767_wire_constant <= "00000001";
    konst_777_wire_constant <= "001";
    konst_785_wire_constant <= "010";
    konst_793_wire_constant <= "011";
    konst_801_wire_constant <= "100";
    konst_807_wire_constant <= "001";
    konst_811_wire_constant <= "00000000000000000000000000000000";
    konst_814_wire_constant <= "010";
    konst_818_wire_constant <= "00000000000000000000000000000000";
    konst_822_wire_constant <= "011";
    konst_826_wire_constant <= "00000000000000000000000000000000";
    konst_829_wire_constant <= "100";
    konst_833_wire_constant <= "00000000000000000000000000000000";
    konst_840_wire_constant <= "001";
    konst_843_wire_constant <= "0";
    konst_846_wire_constant <= "010";
    konst_849_wire_constant <= "0";
    konst_853_wire_constant <= "011";
    konst_856_wire_constant <= "0";
    konst_859_wire_constant <= "100";
    konst_862_wire_constant <= "0";
    konst_872_wire_constant <= "1";
    phi_stmt_657: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_8_659_wire_constant & next_down_counter_772_660_buffered;
      req <= phi_stmt_657_req_0 & phi_stmt_657_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_657",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_657_ack_0,
          idata => idata,
          odata => down_counter_657,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_657
    phi_stmt_661: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_663_wire_constant & RPIPE_noblock_obuf_1_1_665_wire;
      req <= phi_stmt_661_req_0 & phi_stmt_661_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_661",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_661_ack_0,
          idata => idata,
          odata => pkt_1_e_word_661,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_661
    phi_stmt_666: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_668_wire_constant & RPIPE_noblock_obuf_2_1_670_wire;
      req <= phi_stmt_666_req_0 & phi_stmt_666_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_666",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_666_ack_0,
          idata => idata,
          odata => pkt_2_e_word_666,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_666
    phi_stmt_671: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_673_wire_constant & RPIPE_noblock_obuf_3_1_675_wire;
      req <= phi_stmt_671_req_0 & phi_stmt_671_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_671",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_671_ack_0,
          idata => idata,
          odata => pkt_3_e_word_671,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_671
    phi_stmt_676: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_678_wire_constant & RPIPE_noblock_obuf_4_1_680_wire;
      req <= phi_stmt_676_req_0 & phi_stmt_676_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_676",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_676_ack_0,
          idata => idata,
          odata => pkt_4_e_word_676,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_676
    phi_stmt_681: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_3_683_wire_constant & next_active_packet_748_684_buffered;
      req <= phi_stmt_681_req_0 & phi_stmt_681_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_681",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_681_ack_0,
          idata => idata,
          odata => active_packet_681,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_681
    phi_stmt_685: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_3_687_wire_constant & next_pkt_priority_748_688_buffered;
      req <= phi_stmt_685_req_0 & phi_stmt_685_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_685",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_685_ack_0,
          idata => idata,
          odata => pkt_priority_685,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_685
    -- flow-through select operator MUX_716_inst
    MUX_716_wire <= p1_valid_694 when (EQ_u3_u1_713_wire(0) /=  '0') else konst_715_wire_constant;
    -- flow-through select operator MUX_722_inst
    MUX_722_wire <= p2_valid_699 when (EQ_u3_u1_719_wire(0) /=  '0') else konst_721_wire_constant;
    -- flow-through select operator MUX_729_inst
    MUX_729_wire <= p3_valid_704 when (EQ_u3_u1_726_wire(0) /=  '0') else konst_728_wire_constant;
    -- flow-through select operator MUX_735_inst
    MUX_735_wire <= p4_valid_709 when (EQ_u3_u1_732_wire(0) /=  '0') else konst_734_wire_constant;
    -- flow-through select operator MUX_770_inst
    MUX_770_wire <= SUB_u8_u8_768_wire when (valid_active_pkt_word_read_738(0) /=  '0') else down_counter_657;
    -- flow-through select operator MUX_771_inst
    next_down_counter_772 <= konst_764_wire_constant when (started_new_packet_761(0) /=  '0') else MUX_770_wire;
    -- flow-through select operator MUX_812_inst
    MUX_812_wire <= slice_810_wire when (EQ_u3_u1_808_wire(0) /=  '0') else konst_811_wire_constant;
    -- flow-through select operator MUX_819_inst
    MUX_819_wire <= slice_817_wire when (EQ_u3_u1_815_wire(0) /=  '0') else konst_818_wire_constant;
    -- flow-through select operator MUX_827_inst
    MUX_827_wire <= slice_825_wire when (EQ_u3_u1_823_wire(0) /=  '0') else konst_826_wire_constant;
    -- flow-through select operator MUX_834_inst
    MUX_834_wire <= slice_832_wire when (EQ_u3_u1_830_wire(0) /=  '0') else konst_833_wire_constant;
    -- flow-through select operator MUX_844_inst
    MUX_844_wire <= p1_valid_694 when (EQ_u3_u1_841_wire(0) /=  '0') else konst_843_wire_constant;
    -- flow-through select operator MUX_850_inst
    MUX_850_wire <= p2_valid_699 when (EQ_u3_u1_847_wire(0) /=  '0') else konst_849_wire_constant;
    -- flow-through select operator MUX_857_inst
    MUX_857_wire <= p3_valid_704 when (EQ_u3_u1_854_wire(0) /=  '0') else konst_856_wire_constant;
    -- flow-through select operator MUX_863_inst
    MUX_863_wire <= p4_valid_709 when (EQ_u3_u1_860_wire(0) /=  '0') else konst_862_wire_constant;
    -- flow-through slice operator slice_810_inst
    slice_810_wire <= pkt_1_e_word_661(31 downto 0);
    -- flow-through slice operator slice_817_inst
    slice_817_wire <= pkt_2_e_word_666(31 downto 0);
    -- flow-through slice operator slice_825_inst
    slice_825_wire <= pkt_3_e_word_671(31 downto 0);
    -- flow-through slice operator slice_832_inst
    slice_832_wire <= pkt_4_e_word_676(31 downto 0);
    next_active_packet_748_684_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_active_packet_748_684_buf_req_0;
      next_active_packet_748_684_buf_ack_0<= wack(0);
      rreq(0) <= next_active_packet_748_684_buf_req_1;
      next_active_packet_748_684_buf_ack_1<= rack(0);
      next_active_packet_748_684_buf : InterlockBuffer generic map ( -- 
        name => "next_active_packet_748_684_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_active_packet_748,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_active_packet_748_684_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_down_counter_772_660_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_down_counter_772_660_buf_req_0;
      next_down_counter_772_660_buf_ack_0<= wack(0);
      rreq(0) <= next_down_counter_772_660_buf_req_1;
      next_down_counter_772_660_buf_ack_1<= rack(0);
      next_down_counter_772_660_buf : InterlockBuffer generic map ( -- 
        name => "next_down_counter_772_660_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_down_counter_772,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_down_counter_772_660_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_pkt_priority_748_688_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_pkt_priority_748_688_buf_req_0;
      next_pkt_priority_748_688_buf_ack_0<= wack(0);
      rreq(0) <= next_pkt_priority_748_688_buf_req_1;
      next_pkt_priority_748_688_buf_ack_1<= rack(0);
      next_pkt_priority_748_688_buf : InterlockBuffer generic map ( -- 
        name => "next_pkt_priority_748_688_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_pkt_priority_748,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_pkt_priority_748_688_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_655_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_872_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_655_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_655_branch_req_0,
          ack0 => do_while_stmt_655_branch_ack_0,
          ack1 => do_while_stmt_655_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator AND_u1_u1_760_inst
    process(OR_u1_u1_756_wire, EQ_u8_u1_759_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(OR_u1_u1_756_wire, EQ_u8_u1_759_wire, tmp_var);
      started_new_packet_761 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_693_inst
    process(pkt_1_e_word_661) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_1_e_word_661, konst_692_wire_constant, tmp_var);
      p1_valid_694 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_698_inst
    process(pkt_2_e_word_666) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_2_e_word_666, konst_697_wire_constant, tmp_var);
      p2_valid_699 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_703_inst
    process(pkt_3_e_word_671) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_3_e_word_671, konst_702_wire_constant, tmp_var);
      p3_valid_704 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_708_inst
    process(pkt_4_e_word_676) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_4_e_word_676, konst_707_wire_constant, tmp_var);
      p4_valid_709 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_713_inst
    process(active_packet_681) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_681, konst_712_wire_constant, tmp_var);
      EQ_u3_u1_713_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_719_inst
    process(active_packet_681) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_681, konst_718_wire_constant, tmp_var);
      EQ_u3_u1_719_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_726_inst
    process(active_packet_681) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_681, konst_725_wire_constant, tmp_var);
      EQ_u3_u1_726_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_732_inst
    process(active_packet_681) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_681, konst_731_wire_constant, tmp_var);
      EQ_u3_u1_732_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_778_inst
    process(next_active_packet_748) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_748, konst_777_wire_constant, tmp_var);
      EQ_u3_u1_778_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_786_inst
    process(next_active_packet_748) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_748, konst_785_wire_constant, tmp_var);
      EQ_u3_u1_786_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_794_inst
    process(next_active_packet_748) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_748, konst_793_wire_constant, tmp_var);
      EQ_u3_u1_794_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_802_inst
    process(next_active_packet_748) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_748, konst_801_wire_constant, tmp_var);
      EQ_u3_u1_802_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_808_inst
    process(next_active_packet_748) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_748, konst_807_wire_constant, tmp_var);
      EQ_u3_u1_808_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_815_inst
    process(next_active_packet_748) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_748, konst_814_wire_constant, tmp_var);
      EQ_u3_u1_815_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_823_inst
    process(next_active_packet_748) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_748, konst_822_wire_constant, tmp_var);
      EQ_u3_u1_823_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_830_inst
    process(next_active_packet_748) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_748, konst_829_wire_constant, tmp_var);
      EQ_u3_u1_830_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_841_inst
    process(next_active_packet_748) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_748, konst_840_wire_constant, tmp_var);
      EQ_u3_u1_841_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_847_inst
    process(next_active_packet_748) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_748, konst_846_wire_constant, tmp_var);
      EQ_u3_u1_847_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_854_inst
    process(next_active_packet_748) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_748, konst_853_wire_constant, tmp_var);
      EQ_u3_u1_854_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_860_inst
    process(next_active_packet_748) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_748, konst_859_wire_constant, tmp_var);
      EQ_u3_u1_860_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_759_inst
    process(down_counter_657) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(down_counter_657, konst_758_wire_constant, tmp_var);
      EQ_u8_u1_759_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_775_inst
    process(p1_valid_694) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_694, tmp_var);
      NOT_u1_u1_775_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_783_inst
    process(p2_valid_699) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_699, tmp_var);
      NOT_u1_u1_783_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_791_inst
    process(p3_valid_704) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_704, tmp_var);
      NOT_u1_u1_791_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_799_inst
    process(p4_valid_709) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_709, tmp_var);
      NOT_u1_u1_799_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_723_inst
    process(MUX_716_wire, MUX_722_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_716_wire, MUX_722_wire, tmp_var);
      OR_u1_u1_723_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_736_inst
    process(MUX_729_wire, MUX_735_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_729_wire, MUX_735_wire, tmp_var);
      OR_u1_u1_736_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_737_inst
    process(OR_u1_u1_723_wire, OR_u1_u1_736_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_723_wire, OR_u1_u1_736_wire, tmp_var);
      valid_active_pkt_word_read_738 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_752_inst
    process(p1_valid_694, p2_valid_699) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(p1_valid_694, p2_valid_699, tmp_var);
      OR_u1_u1_752_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_755_inst
    process(p3_valid_704, p4_valid_709) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(p3_valid_704, p4_valid_709, tmp_var);
      OR_u1_u1_755_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_756_inst
    process(OR_u1_u1_752_wire, OR_u1_u1_755_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_752_wire, OR_u1_u1_755_wire, tmp_var);
      OR_u1_u1_756_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_779_inst
    process(NOT_u1_u1_775_wire, EQ_u3_u1_778_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_775_wire, EQ_u3_u1_778_wire, tmp_var);
      read_from_1_780 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_787_inst
    process(NOT_u1_u1_783_wire, EQ_u3_u1_786_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_783_wire, EQ_u3_u1_786_wire, tmp_var);
      read_from_2_788 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_795_inst
    process(NOT_u1_u1_791_wire, EQ_u3_u1_794_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_791_wire, EQ_u3_u1_794_wire, tmp_var);
      read_from_3_796 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_803_inst
    process(NOT_u1_u1_799_wire, EQ_u3_u1_802_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_799_wire, EQ_u3_u1_802_wire, tmp_var);
      read_from_4_804 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_851_inst
    process(MUX_844_wire, MUX_850_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_844_wire, MUX_850_wire, tmp_var);
      OR_u1_u1_851_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_864_inst
    process(MUX_857_wire, MUX_863_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_857_wire, MUX_863_wire, tmp_var);
      OR_u1_u1_864_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_865_inst
    process(OR_u1_u1_851_wire, OR_u1_u1_864_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_851_wire, OR_u1_u1_864_wire, tmp_var);
      send_flag_866 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_820_inst
    process(MUX_812_wire, MUX_819_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_812_wire, MUX_819_wire, tmp_var);
      OR_u32_u32_820_wire <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_835_inst
    process(MUX_827_wire, MUX_834_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_827_wire, MUX_834_wire, tmp_var);
      OR_u32_u32_835_wire <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_836_inst
    process(OR_u32_u32_820_wire, OR_u32_u32_835_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u32_u32_820_wire, OR_u32_u32_835_wire, tmp_var);
      data_to_out_837 <= tmp_var; --
    end process;
    -- binary operator SUB_u8_u8_768_inst
    process(down_counter_657) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSub_proc(down_counter_657, konst_767_wire_constant, tmp_var);
      SUB_u8_u8_768_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_noblock_obuf_1_1_665_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_1_1_665_inst_req_0;
      RPIPE_noblock_obuf_1_1_665_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_1_1_665_inst_req_1;
      RPIPE_noblock_obuf_1_1_665_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_1_780(0);
      RPIPE_noblock_obuf_1_1_665_wire <= data_out(32 downto 0);
      noblock_obuf_1_1_read_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_1_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_1_read_0: InputPortRevised -- 
        generic map ( name => "noblock_obuf_1_1_read_0", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_1_1_pipe_read_req(0),
          oack => noblock_obuf_1_1_pipe_read_ack(0),
          odata => noblock_obuf_1_1_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_noblock_obuf_2_1_670_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_2_1_670_inst_req_0;
      RPIPE_noblock_obuf_2_1_670_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_2_1_670_inst_req_1;
      RPIPE_noblock_obuf_2_1_670_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_2_788(0);
      RPIPE_noblock_obuf_2_1_670_wire <= data_out(32 downto 0);
      noblock_obuf_2_1_read_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_1_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_1_read_1: InputPortRevised -- 
        generic map ( name => "noblock_obuf_2_1_read_1", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_2_1_pipe_read_req(0),
          oack => noblock_obuf_2_1_pipe_read_ack(0),
          odata => noblock_obuf_2_1_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_noblock_obuf_3_1_675_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_3_1_675_inst_req_0;
      RPIPE_noblock_obuf_3_1_675_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_3_1_675_inst_req_1;
      RPIPE_noblock_obuf_3_1_675_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_3_796(0);
      RPIPE_noblock_obuf_3_1_675_wire <= data_out(32 downto 0);
      noblock_obuf_3_1_read_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_1_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_1_read_2: InputPortRevised -- 
        generic map ( name => "noblock_obuf_3_1_read_2", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_3_1_pipe_read_req(0),
          oack => noblock_obuf_3_1_pipe_read_ack(0),
          odata => noblock_obuf_3_1_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_noblock_obuf_4_1_680_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_4_1_680_inst_req_0;
      RPIPE_noblock_obuf_4_1_680_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_4_1_680_inst_req_1;
      RPIPE_noblock_obuf_4_1_680_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_4_804(0);
      RPIPE_noblock_obuf_4_1_680_wire <= data_out(32 downto 0);
      noblock_obuf_4_1_read_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_1_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_1_read_3: InputPortRevised -- 
        generic map ( name => "noblock_obuf_4_1_read_3", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_4_1_pipe_read_req(0),
          oack => noblock_obuf_4_1_pipe_read_ack(0),
          odata => noblock_obuf_4_1_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_out_data_1_868_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_out_data_1_868_inst_req_0;
      WPIPE_out_data_1_868_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_out_data_1_868_inst_req_1;
      WPIPE_out_data_1_868_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_flag_866(0);
      data_in <= data_to_out_837;
      out_data_1_write_0_gI: SplitGuardInterface generic map(name => "out_data_1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      out_data_1_write_0: OutputPortRevised -- 
        generic map ( name => "out_data_1", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => out_data_1_pipe_write_req(0),
          oack => out_data_1_pipe_write_ack(0),
          odata => out_data_1_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    volatile_operator_prioritySelect_1970: prioritySelect_Volatile port map(down_counter => down_counter_657, active_packet => active_packet_681, pkt_priority => pkt_priority_685, p1_valid => p1_valid_694, p2_valid => p2_valid_699, p3_valid => p3_valid_704, p4_valid => p4_valid_709, next_active_packet => next_active_packet_748, next_pkt_priority => next_pkt_priority_748); 
    -- 
  end Block; -- data_path
  -- 
end outputPort_1_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity outputPort_2_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    noblock_obuf_1_2_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_2_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_3_2_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_2_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_4_2_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_2_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_2_2_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_2_pipe_read_data : in   std_logic_vector(32 downto 0);
    out_data_2_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_2_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity outputPort_2_Daemon;
architecture outputPort_2_Daemon_arch of outputPort_2_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal outputPort_2_Daemon_CP_1176_start: Boolean;
  signal outputPort_2_Daemon_CP_1176_symbol: Boolean;
  -- volatile/operator module components. 
  component prioritySelect_Volatile is -- 
    port ( -- 
      down_counter : in  std_logic_vector(7 downto 0);
      active_packet : in  std_logic_vector(2 downto 0);
      pkt_priority : in  std_logic_vector(2 downto 0);
      p1_valid : in  std_logic_vector(0 downto 0);
      p2_valid : in  std_logic_vector(0 downto 0);
      p3_valid : in  std_logic_vector(0 downto 0);
      p4_valid : in  std_logic_vector(0 downto 0);
      next_active_packet : out  std_logic_vector(2 downto 0);
      next_pkt_priority : out  std_logic_vector(2 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal phi_stmt_907_req_1 : boolean;
  signal RPIPE_noblock_obuf_1_2_887_inst_ack_1 : boolean;
  signal WPIPE_out_data_2_1090_inst_ack_0 : boolean;
  signal phi_stmt_893_req_1 : boolean;
  signal RPIPE_noblock_obuf_1_2_887_inst_req_1 : boolean;
  signal phi_stmt_893_req_0 : boolean;
  signal phi_stmt_888_req_1 : boolean;
  signal WPIPE_out_data_2_1090_inst_req_0 : boolean;
  signal phi_stmt_893_ack_0 : boolean;
  signal phi_stmt_898_req_1 : boolean;
  signal phi_stmt_903_req_1 : boolean;
  signal phi_stmt_907_ack_0 : boolean;
  signal next_active_packet_970_906_buf_ack_1 : boolean;
  signal RPIPE_noblock_obuf_1_2_887_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_2_887_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_4_2_902_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_2_2_892_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_4_2_902_inst_ack_1 : boolean;
  signal RPIPE_noblock_obuf_2_2_892_inst_ack_1 : boolean;
  signal next_active_packet_970_906_buf_req_1 : boolean;
  signal phi_stmt_888_req_0 : boolean;
  signal phi_stmt_903_req_0 : boolean;
  signal phi_stmt_903_ack_0 : boolean;
  signal phi_stmt_898_req_0 : boolean;
  signal phi_stmt_888_ack_0 : boolean;
  signal WPIPE_out_data_2_1090_inst_req_1 : boolean;
  signal WPIPE_out_data_2_1090_inst_ack_1 : boolean;
  signal next_active_packet_970_906_buf_req_0 : boolean;
  signal next_active_packet_970_906_buf_ack_0 : boolean;
  signal phi_stmt_898_ack_0 : boolean;
  signal phi_stmt_907_req_0 : boolean;
  signal RPIPE_noblock_obuf_3_2_897_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_3_2_897_inst_ack_0 : boolean;
  signal do_while_stmt_877_branch_ack_1 : boolean;
  signal do_while_stmt_877_branch_ack_0 : boolean;
  signal next_pkt_priority_970_910_buf_ack_1 : boolean;
  signal next_pkt_priority_970_910_buf_req_1 : boolean;
  signal RPIPE_noblock_obuf_3_2_897_inst_ack_1 : boolean;
  signal RPIPE_noblock_obuf_3_2_897_inst_req_1 : boolean;
  signal next_pkt_priority_970_910_buf_ack_0 : boolean;
  signal next_pkt_priority_970_910_buf_req_0 : boolean;
  signal RPIPE_noblock_obuf_2_2_892_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_2_2_892_inst_req_0 : boolean;
  signal do_while_stmt_877_branch_req_0 : boolean;
  signal RPIPE_noblock_obuf_4_2_902_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_4_2_902_inst_req_0 : boolean;
  signal phi_stmt_879_req_1 : boolean;
  signal phi_stmt_879_req_0 : boolean;
  signal phi_stmt_879_ack_0 : boolean;
  signal next_down_counter_994_882_buf_req_0 : boolean;
  signal next_down_counter_994_882_buf_ack_0 : boolean;
  signal next_down_counter_994_882_buf_req_1 : boolean;
  signal next_down_counter_994_882_buf_ack_1 : boolean;
  signal phi_stmt_883_req_1 : boolean;
  signal phi_stmt_883_req_0 : boolean;
  signal phi_stmt_883_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "outputPort_2_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  outputPort_2_Daemon_CP_1176_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "outputPort_2_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_2_Daemon_CP_1176_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= outputPort_2_Daemon_CP_1176_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_2_Daemon_CP_1176_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  outputPort_2_Daemon_CP_1176: Block -- control-path 
    signal outputPort_2_Daemon_CP_1176_elements: BooleanArray(161 downto 0);
    -- 
  begin -- 
    outputPort_2_Daemon_CP_1176_elements(0) <= outputPort_2_Daemon_CP_1176_start;
    outputPort_2_Daemon_CP_1176_symbol <= outputPort_2_Daemon_CP_1176_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_876/$entry
      -- CP-element group 0: 	 branch_block_stmt_876/branch_block_stmt_876__entry__
      -- CP-element group 0: 	 branch_block_stmt_876/do_while_stmt_877__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	161 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_876/$exit
      -- CP-element group 1: 	 branch_block_stmt_876/branch_block_stmt_876__exit__
      -- CP-element group 1: 	 branch_block_stmt_876/do_while_stmt_877__exit__
      -- 
    outputPort_2_Daemon_CP_1176_elements(1) <= outputPort_2_Daemon_CP_1176_elements(161);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_876/do_while_stmt_877/$entry
      -- CP-element group 2: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877__entry__
      -- 
    outputPort_2_Daemon_CP_1176_elements(2) <= outputPort_2_Daemon_CP_1176_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	161 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877__exit__
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_876/do_while_stmt_877/loop_back
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	159 
    -- CP-element group 5: 	160 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_876/do_while_stmt_877/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_876/do_while_stmt_877/condition_done
      -- CP-element group 5: 	 branch_block_stmt_876/do_while_stmt_877/loop_taken/$entry
      -- 
    outputPort_2_Daemon_CP_1176_elements(5) <= outputPort_2_Daemon_CP_1176_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	158 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_876/do_while_stmt_877/loop_body_done
      -- 
    outputPort_2_Daemon_CP_1176_elements(6) <= outputPort_2_Daemon_CP_1176_elements(158);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	141 
    -- CP-element group 7: 	103 
    -- CP-element group 7: 	124 
    -- CP-element group 7: 	21 
    -- CP-element group 7: 	40 
    -- CP-element group 7: 	82 
    -- CP-element group 7: 	61 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/back_edge_to_loop_body
      -- 
    outputPort_2_Daemon_CP_1176_elements(7) <= outputPort_2_Daemon_CP_1176_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	143 
    -- CP-element group 8: 	84 
    -- CP-element group 8: 	23 
    -- CP-element group 8: 	42 
    -- CP-element group 8: 	126 
    -- CP-element group 8: 	105 
    -- CP-element group 8: 	63 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/first_time_through_loop_body
      -- 
    outputPort_2_Daemon_CP_1176_elements(8) <= outputPort_2_Daemon_CP_1176_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	157 
    -- CP-element group 9: 	97 
    -- CP-element group 9: 	77 
    -- CP-element group 9: 	76 
    -- CP-element group 9: 	119 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	34 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	118 
    -- CP-element group 9: 	137 
    -- CP-element group 9: 	138 
    -- CP-element group 9: 	98 
    -- CP-element group 9: 	55 
    -- CP-element group 9: 	56 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/loop_body_start
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	157 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/condition_evaluated
      -- 
    condition_evaluated_1200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(10), ack => do_while_stmt_877_branch_req_0); -- 
    outputPort_2_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(157) & outputPort_2_Daemon_CP_1176_elements(14);
      gj_outputPort_2_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	97 
    -- CP-element group 11: 	76 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	118 
    -- CP-element group 11: 	137 
    -- CP-element group 11: 	55 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	99 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	120 
    -- CP-element group 11: 	78 
    -- CP-element group 11: 	57 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_907_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/aggregated_phi_sample_req
      -- 
    outputPort_2_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(97) & outputPort_2_Daemon_CP_1176_elements(76) & outputPort_2_Daemon_CP_1176_elements(15) & outputPort_2_Daemon_CP_1176_elements(34) & outputPort_2_Daemon_CP_1176_elements(118) & outputPort_2_Daemon_CP_1176_elements(137) & outputPort_2_Daemon_CP_1176_elements(55) & outputPort_2_Daemon_CP_1176_elements(14);
      gj_outputPort_2_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	139 
    -- CP-element group 12: 	100 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	37 
    -- CP-element group 12: 	121 
    -- CP-element group 12: 	79 
    -- CP-element group 12: 	58 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	158 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	97 
    -- CP-element group 12: 	76 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	34 
    -- CP-element group 12: 	118 
    -- CP-element group 12: 	137 
    -- CP-element group 12: 	55 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_888_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_903_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_893_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_907_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_898_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_879_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_883_sample_completed_
      -- 
    outputPort_2_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(139) & outputPort_2_Daemon_CP_1176_elements(100) & outputPort_2_Daemon_CP_1176_elements(18) & outputPort_2_Daemon_CP_1176_elements(37) & outputPort_2_Daemon_CP_1176_elements(121) & outputPort_2_Daemon_CP_1176_elements(79) & outputPort_2_Daemon_CP_1176_elements(58);
      gj_outputPort_2_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	77 
    -- CP-element group 13: 	119 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	35 
    -- CP-element group 13: 	138 
    -- CP-element group 13: 	98 
    -- CP-element group 13: 	56 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	101 
    -- CP-element group 13: 	19 
    -- CP-element group 13: 	38 
    -- CP-element group 13: 	122 
    -- CP-element group 13: 	80 
    -- CP-element group 13: 	59 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_907_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/aggregated_phi_update_req
      -- 
    outputPort_2_Daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(77) & outputPort_2_Daemon_CP_1176_elements(119) & outputPort_2_Daemon_CP_1176_elements(16) & outputPort_2_Daemon_CP_1176_elements(35) & outputPort_2_Daemon_CP_1176_elements(138) & outputPort_2_Daemon_CP_1176_elements(98) & outputPort_2_Daemon_CP_1176_elements(56);
      gj_outputPort_2_Daemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	140 
    -- CP-element group 14: 	102 
    -- CP-element group 14: 	123 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	81 
    -- CP-element group 14: 	60 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/aggregated_phi_update_ack
      -- 
    outputPort_2_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(140) & outputPort_2_Daemon_CP_1176_elements(102) & outputPort_2_Daemon_CP_1176_elements(123) & outputPort_2_Daemon_CP_1176_elements(20) & outputPort_2_Daemon_CP_1176_elements(39) & outputPort_2_Daemon_CP_1176_elements(81) & outputPort_2_Daemon_CP_1176_elements(60);
      gj_outputPort_2_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_879_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	155 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_879_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(155);
      gj_outputPort_2_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_879_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(17) <= outputPort_2_Daemon_CP_1176_elements(11);
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_879_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_879_update_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(19) <= outputPort_2_Daemon_CP_1176_elements(13);
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	154 
    -- CP-element group 20: 	14 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_879_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_879_update_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_879_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(21) <= outputPort_2_Daemon_CP_1176_elements(7);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_879_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_879_loopback_sample_req_ps
      -- 
    phi_stmt_879_loopback_sample_req_1215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_879_loopback_sample_req_1215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(22), ack => phi_stmt_879_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_879_entry_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(23) <= outputPort_2_Daemon_CP_1176_elements(8);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_879_entry_sample_req
      -- CP-element group 24: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_879_entry_sample_req_ps
      -- 
    phi_stmt_879_entry_sample_req_1218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_879_entry_sample_req_1218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(24), ack => phi_stmt_879_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_879_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_879_phi_mux_ack_ps
      -- 
    phi_stmt_879_phi_mux_ack_1221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_879_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_8_881_sample_start__ps
      -- CP-element group 26: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_8_881_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_8_881_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_8_881_sample_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_8_881_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_8_881_update_start_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_8_881_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(28) <= outputPort_2_Daemon_CP_1176_elements(29);
    -- CP-element group 29:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	28 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_8_881_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(29) is a control-delay.
    cp_element_29_delay: control_delay_element  generic map(name => " 29_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_1176_elements(27), ack => outputPort_2_Daemon_CP_1176_elements(29), clk => clk, reset =>reset);
    -- CP-element group 30:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_down_counter_882_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_down_counter_882_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_down_counter_882_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_down_counter_882_Sample/req
      -- 
    req_1242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(30), ack => next_down_counter_994_882_buf_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_down_counter_882_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_down_counter_882_update_start_
      -- CP-element group 31: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_down_counter_882_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_down_counter_882_Update/req
      -- 
    req_1247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(31), ack => next_down_counter_994_882_buf_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_down_counter_882_sample_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_down_counter_882_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_down_counter_882_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_down_counter_882_Sample/ack
      -- 
    ack_1243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_994_882_buf_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(32)); -- 
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_down_counter_882_update_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_down_counter_882_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_down_counter_882_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_down_counter_882_Update/ack
      -- 
    ack_1248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_994_882_buf_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(33)); -- 
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	9 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	12 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	11 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_883_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	155 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	13 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_883_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(155);
      gj_outputPort_2_Daemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	11 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_883_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(36) <= outputPort_2_Daemon_CP_1176_elements(11);
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	12 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_883_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_883_update_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(38) <= outputPort_2_Daemon_CP_1176_elements(13);
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	154 
    -- CP-element group 39: 	14 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_883_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_883_update_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	7 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_883_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(40) <= outputPort_2_Daemon_CP_1176_elements(7);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_883_loopback_sample_req
      -- CP-element group 41: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_883_loopback_sample_req_ps
      -- 
    phi_stmt_883_loopback_sample_req_1259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_883_loopback_sample_req_1259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(41), ack => phi_stmt_883_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	8 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_883_entry_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(42) <= outputPort_2_Daemon_CP_1176_elements(8);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_883_entry_sample_req
      -- CP-element group 43: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_883_entry_sample_req_ps
      -- 
    phi_stmt_883_entry_sample_req_1262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_883_entry_sample_req_1262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(43), ack => phi_stmt_883_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_883_phi_mux_ack
      -- CP-element group 44: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_883_phi_mux_ack_ps
      -- 
    phi_stmt_883_phi_mux_ack_1265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_883_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_885_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_885_sample_start__ps
      -- CP-element group 45: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_885_sample_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_885_sample_start_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_885_update_start_
      -- CP-element group 46: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_885_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_885_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(47) <= outputPort_2_Daemon_CP_1176_elements(48);
    -- CP-element group 48:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	47 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_885_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(48) is a control-delay.
    cp_element_48_delay: control_delay_element  generic map(name => " 48_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_1176_elements(46), ack => outputPort_2_Daemon_CP_1176_elements(48), clk => clk, reset =>reset);
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_1_2_887_sample_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_1_2_887_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	54 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_1_2_887_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_1_2_887_Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_1_2_887_Sample/$entry
      -- 
    rr_1286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(51), ack => RPIPE_noblock_obuf_1_2_887_inst_req_0); -- 
    outputPort_2_Daemon_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(49) & outputPort_2_Daemon_CP_1176_elements(54);
      gj_outputPort_2_Daemon_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: 	53 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_1_2_887_update_start_
      -- CP-element group 52: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_1_2_887_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_1_2_887_Update/$entry
      -- 
    cr_1291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(52), ack => RPIPE_noblock_obuf_1_2_887_inst_req_1); -- 
    outputPort_2_Daemon_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(50) & outputPort_2_Daemon_CP_1176_elements(53);
      gj_outputPort_2_Daemon_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	52 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_1_2_887_sample_completed__ps
      -- CP-element group 53: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_1_2_887_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_1_2_887_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_1_2_887_sample_completed_
      -- 
    ra_1287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_2_887_inst_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(53)); -- 
    -- CP-element group 54:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	51 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_1_2_887_update_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_1_2_887_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_1_2_887_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_1_2_887_update_completed_
      -- 
    ca_1292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_2_887_inst_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(54)); -- 
    -- CP-element group 55:  join  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	9 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	12 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	11 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_888_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	9 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	155 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	13 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_888_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(155);
      gj_outputPort_2_Daemon_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	11 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_888_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(57) <= outputPort_2_Daemon_CP_1176_elements(11);
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	12 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_888_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	13 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_888_update_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(59) <= outputPort_2_Daemon_CP_1176_elements(13);
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	154 
    -- CP-element group 60: 	14 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_888_update_completed__ps
      -- CP-element group 60: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_888_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	7 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_888_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(61) <= outputPort_2_Daemon_CP_1176_elements(7);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_888_loopback_sample_req_ps
      -- CP-element group 62: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_888_loopback_sample_req
      -- 
    phi_stmt_888_loopback_sample_req_1303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_888_loopback_sample_req_1303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(62), ack => phi_stmt_888_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	8 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_888_entry_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(63) <= outputPort_2_Daemon_CP_1176_elements(8);
    -- CP-element group 64:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_888_entry_sample_req
      -- CP-element group 64: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_888_entry_sample_req_ps
      -- 
    phi_stmt_888_entry_sample_req_1306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_888_entry_sample_req_1306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(64), ack => phi_stmt_888_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_888_phi_mux_ack
      -- CP-element group 65: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_888_phi_mux_ack_ps
      -- 
    phi_stmt_888_phi_mux_ack_1309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_888_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(65)); -- 
    -- CP-element group 66:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_890_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_890_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_890_sample_start__ps
      -- CP-element group 66: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_890_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_890_update_start_
      -- CP-element group 67: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_890_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_890_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(68) <= outputPort_2_Daemon_CP_1176_elements(69);
    -- CP-element group 69:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	68 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_890_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(69) is a control-delay.
    cp_element_69_delay: control_delay_element  generic map(name => " 69_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_1176_elements(67), ack => outputPort_2_Daemon_CP_1176_elements(69), clk => clk, reset =>reset);
    -- CP-element group 70:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_2_2_892_sample_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(70) is bound as output of CP function.
    -- CP-element group 71:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_2_2_892_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: marked-predecessors 
    -- CP-element group 72: 	75 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_2_2_892_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_2_2_892_Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_2_2_892_Sample/$entry
      -- 
    rr_1330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(72), ack => RPIPE_noblock_obuf_2_2_892_inst_req_0); -- 
    outputPort_2_Daemon_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(70) & outputPort_2_Daemon_CP_1176_elements(75);
      gj_outputPort_2_Daemon_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: 	74 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_2_2_892_update_start_
      -- CP-element group 73: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_2_2_892_Update/cr
      -- CP-element group 73: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_2_2_892_Update/$entry
      -- 
    cr_1335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(73), ack => RPIPE_noblock_obuf_2_2_892_inst_req_1); -- 
    outputPort_2_Daemon_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(71) & outputPort_2_Daemon_CP_1176_elements(74);
      gj_outputPort_2_Daemon_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	73 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_2_2_892_sample_completed__ps
      -- CP-element group 74: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_2_2_892_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_2_2_892_Sample/ra
      -- CP-element group 74: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_2_2_892_Sample/$exit
      -- 
    ra_1331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_2_892_inst_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(74)); -- 
    -- CP-element group 75:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	72 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_2_2_892_update_completed__ps
      -- CP-element group 75: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_2_2_892_Update/ca
      -- CP-element group 75: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_2_2_892_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_2_2_892_update_completed_
      -- 
    ca_1336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_2_892_inst_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(75)); -- 
    -- CP-element group 76:  join  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	9 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	12 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	11 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_893_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	9 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	155 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	13 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_893_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(155);
      gj_outputPort_2_Daemon_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	11 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_893_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(78) <= outputPort_2_Daemon_CP_1176_elements(11);
    -- CP-element group 79:  join  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	12 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_893_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	13 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_893_update_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(80) <= outputPort_2_Daemon_CP_1176_elements(13);
    -- CP-element group 81:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	154 
    -- CP-element group 81: 	14 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_893_update_completed__ps
      -- CP-element group 81: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_893_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	7 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_893_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(82) <= outputPort_2_Daemon_CP_1176_elements(7);
    -- CP-element group 83:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_893_loopback_sample_req_ps
      -- CP-element group 83: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_893_loopback_sample_req
      -- 
    phi_stmt_893_loopback_sample_req_1347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_893_loopback_sample_req_1347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(83), ack => phi_stmt_893_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(83) is bound as output of CP function.
    -- CP-element group 84:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	8 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_893_entry_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(84) <= outputPort_2_Daemon_CP_1176_elements(8);
    -- CP-element group 85:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_893_entry_sample_req_ps
      -- CP-element group 85: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_893_entry_sample_req
      -- 
    phi_stmt_893_entry_sample_req_1350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_893_entry_sample_req_1350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(85), ack => phi_stmt_893_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_893_phi_mux_ack_ps
      -- CP-element group 86: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_893_phi_mux_ack
      -- 
    phi_stmt_893_phi_mux_ack_1353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_893_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(86)); -- 
    -- CP-element group 87:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_895_sample_completed__ps
      -- CP-element group 87: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_895_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_895_sample_start__ps
      -- CP-element group 87: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_895_sample_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_895_update_start__ps
      -- CP-element group 88: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_895_update_start_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	90 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_895_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(89) <= outputPort_2_Daemon_CP_1176_elements(90);
    -- CP-element group 90:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	89 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_895_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(90) is a control-delay.
    cp_element_90_delay: control_delay_element  generic map(name => " 90_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_1176_elements(88), ack => outputPort_2_Daemon_CP_1176_elements(90), clk => clk, reset =>reset);
    -- CP-element group 91:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_3_2_897_sample_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(91) is bound as output of CP function.
    -- CP-element group 92:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_3_2_897_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(92) is bound as output of CP function.
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	96 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_3_2_897_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_3_2_897_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_3_2_897_Sample/rr
      -- 
    rr_1374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(93), ack => RPIPE_noblock_obuf_3_2_897_inst_req_0); -- 
    outputPort_2_Daemon_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(91) & outputPort_2_Daemon_CP_1176_elements(96);
      gj_outputPort_2_Daemon_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	95 
    -- CP-element group 94: 	92 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_3_2_897_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_3_2_897_update_start_
      -- CP-element group 94: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_3_2_897_Update/cr
      -- 
    cr_1379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(94), ack => RPIPE_noblock_obuf_3_2_897_inst_req_1); -- 
    outputPort_2_Daemon_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(95) & outputPort_2_Daemon_CP_1176_elements(92);
      gj_outputPort_2_Daemon_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	94 
    -- CP-element group 95:  members (4) 
      -- CP-element group 95: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_3_2_897_sample_completed__ps
      -- CP-element group 95: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_3_2_897_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_3_2_897_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_3_2_897_Sample/ra
      -- 
    ra_1375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_2_897_inst_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(95)); -- 
    -- CP-element group 96:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	93 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_3_2_897_update_completed__ps
      -- CP-element group 96: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_3_2_897_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_3_2_897_Update/ca
      -- CP-element group 96: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_3_2_897_Update/$exit
      -- 
    ca_1380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_2_897_inst_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(96)); -- 
    -- CP-element group 97:  join  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	9 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	12 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	11 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_898_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	9 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	155 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	13 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_898_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_2_Daemon_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(155);
      gj_outputPort_2_Daemon_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	11 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_898_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(99) <= outputPort_2_Daemon_CP_1176_elements(11);
    -- CP-element group 100:  join  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	12 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_898_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(100) is bound as output of CP function.
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	13 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_898_update_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(101) <= outputPort_2_Daemon_CP_1176_elements(13);
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	154 
    -- CP-element group 102: 	14 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_898_update_completed__ps
      -- CP-element group 102: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_898_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(102) is bound as output of CP function.
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	7 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_898_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(103) <= outputPort_2_Daemon_CP_1176_elements(7);
    -- CP-element group 104:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_898_loopback_sample_req_ps
      -- CP-element group 104: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_898_loopback_sample_req
      -- 
    phi_stmt_898_loopback_sample_req_1391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_898_loopback_sample_req_1391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(104), ack => phi_stmt_898_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(104) is bound as output of CP function.
    -- CP-element group 105:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	8 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_898_entry_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(105) <= outputPort_2_Daemon_CP_1176_elements(8);
    -- CP-element group 106:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_898_entry_sample_req
      -- CP-element group 106: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_898_entry_sample_req_ps
      -- 
    phi_stmt_898_entry_sample_req_1394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_898_entry_sample_req_1394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(106), ack => phi_stmt_898_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_898_phi_mux_ack
      -- CP-element group 107: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_898_phi_mux_ack_ps
      -- 
    phi_stmt_898_phi_mux_ack_1397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_898_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(107)); -- 
    -- CP-element group 108:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_900_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_900_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_900_sample_completed__ps
      -- CP-element group 108: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_900_sample_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(108) is bound as output of CP function.
    -- CP-element group 109:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_900_update_start_
      -- CP-element group 109: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_900_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	111 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_900_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(110) <= outputPort_2_Daemon_CP_1176_elements(111);
    -- CP-element group 111:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	110 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_33_900_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(111) is a control-delay.
    cp_element_111_delay: control_delay_element  generic map(name => " 111_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_1176_elements(109), ack => outputPort_2_Daemon_CP_1176_elements(111), clk => clk, reset =>reset);
    -- CP-element group 112:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_4_2_902_sample_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(112) is bound as output of CP function.
    -- CP-element group 113:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_4_2_902_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(113) is bound as output of CP function.
    -- CP-element group 114:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: marked-predecessors 
    -- CP-element group 114: 	117 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_4_2_902_Sample/rr
      -- CP-element group 114: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_4_2_902_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_4_2_902_sample_start_
      -- 
    rr_1418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(114), ack => RPIPE_noblock_obuf_4_2_902_inst_req_0); -- 
    outputPort_2_Daemon_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(112) & outputPort_2_Daemon_CP_1176_elements(117);
      gj_outputPort_2_Daemon_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	116 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_4_2_902_Update/cr
      -- CP-element group 115: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_4_2_902_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_4_2_902_update_start_
      -- 
    cr_1423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(115), ack => RPIPE_noblock_obuf_4_2_902_inst_req_1); -- 
    outputPort_2_Daemon_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(113) & outputPort_2_Daemon_CP_1176_elements(116);
      gj_outputPort_2_Daemon_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	115 
    -- CP-element group 116:  members (4) 
      -- CP-element group 116: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_4_2_902_Sample/ra
      -- CP-element group 116: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_4_2_902_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_4_2_902_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_4_2_902_sample_completed__ps
      -- 
    ra_1419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_2_902_inst_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(116)); -- 
    -- CP-element group 117:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: marked-successors 
    -- CP-element group 117: 	114 
    -- CP-element group 117:  members (4) 
      -- CP-element group 117: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_4_2_902_Update/ca
      -- CP-element group 117: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_4_2_902_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_4_2_902_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/RPIPE_noblock_obuf_4_2_902_update_completed__ps
      -- 
    ca_1424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_2_902_inst_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(117)); -- 
    -- CP-element group 118:  join  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	9 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	12 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	11 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_903_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  join  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	9 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	155 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	13 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_903_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(155);
      gj_outputPort_2_Daemon_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	11 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_903_sample_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(120) <= outputPort_2_Daemon_CP_1176_elements(11);
    -- CP-element group 121:  join  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	12 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_903_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(121) is bound as output of CP function.
    -- CP-element group 122:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	13 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_903_update_start__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(122) <= outputPort_2_Daemon_CP_1176_elements(13);
    -- CP-element group 123:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	154 
    -- CP-element group 123: 	14 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_903_update_completed__ps
      -- CP-element group 123: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_903_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(123) is bound as output of CP function.
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	7 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_903_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(124) <= outputPort_2_Daemon_CP_1176_elements(7);
    -- CP-element group 125:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_903_loopback_sample_req_ps
      -- CP-element group 125: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_903_loopback_sample_req
      -- 
    phi_stmt_903_loopback_sample_req_1435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_903_loopback_sample_req_1435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(125), ack => phi_stmt_903_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(125) is bound as output of CP function.
    -- CP-element group 126:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	8 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_903_entry_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(126) <= outputPort_2_Daemon_CP_1176_elements(8);
    -- CP-element group 127:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_903_entry_sample_req
      -- CP-element group 127: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_903_entry_sample_req_ps
      -- 
    phi_stmt_903_entry_sample_req_1438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_903_entry_sample_req_1438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(127), ack => phi_stmt_903_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(127) is bound as output of CP function.
    -- CP-element group 128:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_903_phi_mux_ack
      -- CP-element group 128: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_903_phi_mux_ack_ps
      -- 
    phi_stmt_903_phi_mux_ack_1441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_903_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(128)); -- 
    -- CP-element group 129:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (4) 
      -- CP-element group 129: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_3_905_sample_start__ps
      -- CP-element group 129: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_3_905_sample_completed__ps
      -- CP-element group 129: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_3_905_sample_start_
      -- CP-element group 129: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_3_905_sample_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(129) is bound as output of CP function.
    -- CP-element group 130:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (2) 
      -- CP-element group 130: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_3_905_update_start__ps
      -- CP-element group 130: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_3_905_update_start_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(130) is bound as output of CP function.
    -- CP-element group 131:  join  transition  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	132 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_3_905_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(131) <= outputPort_2_Daemon_CP_1176_elements(132);
    -- CP-element group 132:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	131 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_3_905_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(132) is a control-delay.
    cp_element_132_delay: control_delay_element  generic map(name => " 132_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_1176_elements(130), ack => outputPort_2_Daemon_CP_1176_elements(132), clk => clk, reset =>reset);
    -- CP-element group 133:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	135 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_active_packet_906_sample_start__ps
      -- CP-element group 133: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_active_packet_906_sample_start_
      -- CP-element group 133: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_active_packet_906_Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_active_packet_906_Sample/req
      -- 
    req_1462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(133), ack => next_active_packet_970_906_buf_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(133) is bound as output of CP function.
    -- CP-element group 134:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_active_packet_906_Update/req
      -- CP-element group 134: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_active_packet_906_update_start__ps
      -- CP-element group 134: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_active_packet_906_update_start_
      -- CP-element group 134: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_active_packet_906_Update/$entry
      -- 
    req_1467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(134), ack => next_active_packet_970_906_buf_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(134) is bound as output of CP function.
    -- CP-element group 135:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	133 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (4) 
      -- CP-element group 135: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_active_packet_906_sample_completed__ps
      -- CP-element group 135: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_active_packet_906_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_active_packet_906_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_active_packet_906_Sample/ack
      -- 
    ack_1463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_970_906_buf_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(135)); -- 
    -- CP-element group 136:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (4) 
      -- CP-element group 136: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_active_packet_906_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_active_packet_906_Update/ack
      -- CP-element group 136: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_active_packet_906_update_completed__ps
      -- CP-element group 136: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_active_packet_906_update_completed_
      -- 
    ack_1468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_970_906_buf_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(136)); -- 
    -- CP-element group 137:  join  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	9 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	12 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	11 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_907_sample_start_
      -- 
    outputPort_2_Daemon_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(12);
      gj_outputPort_2_Daemon_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  join  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	9 
    -- CP-element group 138: marked-predecessors 
    -- CP-element group 138: 	155 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	13 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_907_update_start_
      -- 
    outputPort_2_Daemon_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(9) & outputPort_2_Daemon_CP_1176_elements(155);
      gj_outputPort_2_Daemon_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 139:  join  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	12 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_907_sample_completed__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(139) is bound as output of CP function.
    -- CP-element group 140:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	154 
    -- CP-element group 140: 	14 
    -- CP-element group 140:  members (2) 
      -- CP-element group 140: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_907_update_completed__ps
      -- CP-element group 140: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_907_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(140) is bound as output of CP function.
    -- CP-element group 141:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	7 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_907_loopback_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(141) <= outputPort_2_Daemon_CP_1176_elements(7);
    -- CP-element group 142:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_907_loopback_sample_req
      -- CP-element group 142: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_907_loopback_sample_req_ps
      -- 
    phi_stmt_907_loopback_sample_req_1479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_907_loopback_sample_req_1479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(142), ack => phi_stmt_907_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(142) is bound as output of CP function.
    -- CP-element group 143:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	8 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_907_entry_trigger
      -- 
    outputPort_2_Daemon_CP_1176_elements(143) <= outputPort_2_Daemon_CP_1176_elements(8);
    -- CP-element group 144:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_907_entry_sample_req
      -- CP-element group 144: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_907_entry_sample_req_ps
      -- 
    phi_stmt_907_entry_sample_req_1482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_907_entry_sample_req_1482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(144), ack => phi_stmt_907_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_907_phi_mux_ack
      -- CP-element group 145: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/phi_stmt_907_phi_mux_ack_ps
      -- 
    phi_stmt_907_phi_mux_ack_1485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_907_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(145)); -- 
    -- CP-element group 146:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (4) 
      -- CP-element group 146: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_3_909_sample_completed_
      -- CP-element group 146: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_3_909_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_3_909_sample_completed__ps
      -- CP-element group 146: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_3_909_sample_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(146) is bound as output of CP function.
    -- CP-element group 147:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (2) 
      -- CP-element group 147: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_3_909_update_start_
      -- CP-element group 147: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_3_909_update_start__ps
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(147) is bound as output of CP function.
    -- CP-element group 148:  join  transition  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	149 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (1) 
      -- CP-element group 148: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_3_909_update_completed__ps
      -- 
    outputPort_2_Daemon_CP_1176_elements(148) <= outputPort_2_Daemon_CP_1176_elements(149);
    -- CP-element group 149:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	148 
    -- CP-element group 149:  members (1) 
      -- CP-element group 149: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_ZERO_3_909_update_completed_
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(149) is a control-delay.
    cp_element_149_delay: control_delay_element  generic map(name => " 149_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_1176_elements(147), ack => outputPort_2_Daemon_CP_1176_elements(149), clk => clk, reset =>reset);
    -- CP-element group 150:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (4) 
      -- CP-element group 150: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_pkt_priority_910_sample_start__ps
      -- CP-element group 150: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_pkt_priority_910_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_pkt_priority_910_Sample/req
      -- CP-element group 150: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_pkt_priority_910_Sample/$entry
      -- 
    req_1506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(150), ack => next_pkt_priority_970_910_buf_req_0); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(150) is bound as output of CP function.
    -- CP-element group 151:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (4) 
      -- CP-element group 151: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_pkt_priority_910_update_start__ps
      -- CP-element group 151: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_pkt_priority_910_update_start_
      -- CP-element group 151: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_pkt_priority_910_Update/req
      -- CP-element group 151: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_pkt_priority_910_Update/$entry
      -- 
    req_1511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(151), ack => next_pkt_priority_970_910_buf_req_1); -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(151) is bound as output of CP function.
    -- CP-element group 152:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (4) 
      -- CP-element group 152: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_pkt_priority_910_sample_completed__ps
      -- CP-element group 152: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_pkt_priority_910_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_pkt_priority_910_Sample/ack
      -- CP-element group 152: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_pkt_priority_910_Sample/$exit
      -- 
    ack_1507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pkt_priority_970_910_buf_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(152)); -- 
    -- CP-element group 153:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (4) 
      -- CP-element group 153: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_pkt_priority_910_update_completed__ps
      -- CP-element group 153: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_pkt_priority_910_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_pkt_priority_910_Update/ack
      -- CP-element group 153: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/R_next_pkt_priority_910_Update/$exit
      -- 
    ack_1512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pkt_priority_970_910_buf_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	140 
    -- CP-element group 154: 	102 
    -- CP-element group 154: 	123 
    -- CP-element group 154: 	20 
    -- CP-element group 154: 	39 
    -- CP-element group 154: 	81 
    -- CP-element group 154: 	60 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/WPIPE_out_data_2_1090_Sample/req
      -- CP-element group 154: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/WPIPE_out_data_2_1090_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/WPIPE_out_data_2_1090_sample_start_
      -- 
    req_1521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(154), ack => WPIPE_out_data_2_1090_inst_req_0); -- 
    outputPort_2_Daemon_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(140) & outputPort_2_Daemon_CP_1176_elements(102) & outputPort_2_Daemon_CP_1176_elements(123) & outputPort_2_Daemon_CP_1176_elements(20) & outputPort_2_Daemon_CP_1176_elements(39) & outputPort_2_Daemon_CP_1176_elements(81) & outputPort_2_Daemon_CP_1176_elements(60) & outputPort_2_Daemon_CP_1176_elements(156);
      gj_outputPort_2_Daemon_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	77 
    -- CP-element group 155: 	119 
    -- CP-element group 155: 	16 
    -- CP-element group 155: 	35 
    -- CP-element group 155: 	138 
    -- CP-element group 155: 	98 
    -- CP-element group 155: 	56 
    -- CP-element group 155:  members (6) 
      -- CP-element group 155: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/WPIPE_out_data_2_1090_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/WPIPE_out_data_2_1090_Sample/ack
      -- CP-element group 155: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/WPIPE_out_data_2_1090_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/WPIPE_out_data_2_1090_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/WPIPE_out_data_2_1090_update_start_
      -- CP-element group 155: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/WPIPE_out_data_2_1090_Update/req
      -- 
    ack_1522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_2_1090_inst_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(155)); -- 
    req_1526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_2_Daemon_CP_1176_elements(155), ack => WPIPE_out_data_2_1090_inst_req_1); -- 
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	154 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/WPIPE_out_data_2_1090_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/WPIPE_out_data_2_1090_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/WPIPE_out_data_2_1090_Update/ack
      -- 
    ack_1527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_2_1090_inst_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(156)); -- 
    -- CP-element group 157:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	9 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	10 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group outputPort_2_Daemon_CP_1176_elements(157) is a control-delay.
    cp_element_157_delay: control_delay_element  generic map(name => " 157_delay", delay_value => 1)  port map(req => outputPort_2_Daemon_CP_1176_elements(9), ack => outputPort_2_Daemon_CP_1176_elements(157), clk => clk, reset =>reset);
    -- CP-element group 158:  join  transition  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	12 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	6 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_876/do_while_stmt_877/do_while_stmt_877_loop_body/$exit
      -- 
    outputPort_2_Daemon_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_2_Daemon_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_2_Daemon_CP_1176_elements(12) & outputPort_2_Daemon_CP_1176_elements(156);
      gj_outputPort_2_Daemon_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	5 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (2) 
      -- CP-element group 159: 	 branch_block_stmt_876/do_while_stmt_877/loop_exit/ack
      -- CP-element group 159: 	 branch_block_stmt_876/do_while_stmt_877/loop_exit/$exit
      -- 
    ack_1532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_877_branch_ack_0, ack => outputPort_2_Daemon_CP_1176_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	5 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (2) 
      -- CP-element group 160: 	 branch_block_stmt_876/do_while_stmt_877/loop_taken/ack
      -- CP-element group 160: 	 branch_block_stmt_876/do_while_stmt_877/loop_taken/$exit
      -- 
    ack_1536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_877_branch_ack_1, ack => outputPort_2_Daemon_CP_1176_elements(160)); -- 
    -- CP-element group 161:  transition  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	3 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	1 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_876/do_while_stmt_877/$exit
      -- 
    outputPort_2_Daemon_CP_1176_elements(161) <= outputPort_2_Daemon_CP_1176_elements(3);
    outputPort_2_Daemon_do_while_stmt_877_terminator_1537: loop_terminator -- 
      generic map (name => " outputPort_2_Daemon_do_while_stmt_877_terminator_1537", max_iterations_in_flight =>7) 
      port map(loop_body_exit => outputPort_2_Daemon_CP_1176_elements(6),loop_continue => outputPort_2_Daemon_CP_1176_elements(160),loop_terminate => outputPort_2_Daemon_CP_1176_elements(159),loop_back => outputPort_2_Daemon_CP_1176_elements(4),loop_exit => outputPort_2_Daemon_CP_1176_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_879_phi_seq_1249_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_1176_elements(23);
      outputPort_2_Daemon_CP_1176_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(26);
      outputPort_2_Daemon_CP_1176_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(28);
      outputPort_2_Daemon_CP_1176_elements(24) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_1176_elements(21);
      outputPort_2_Daemon_CP_1176_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(32);
      outputPort_2_Daemon_CP_1176_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(33);
      outputPort_2_Daemon_CP_1176_elements(22) <= phi_mux_reqs(1);
      phi_stmt_879_phi_seq_1249 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_879_phi_seq_1249") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_1176_elements(17), 
          phi_sample_ack => outputPort_2_Daemon_CP_1176_elements(18), 
          phi_update_req => outputPort_2_Daemon_CP_1176_elements(19), 
          phi_update_ack => outputPort_2_Daemon_CP_1176_elements(20), 
          phi_mux_ack => outputPort_2_Daemon_CP_1176_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_883_phi_seq_1293_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_1176_elements(42);
      outputPort_2_Daemon_CP_1176_elements(45)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(45);
      outputPort_2_Daemon_CP_1176_elements(46)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(47);
      outputPort_2_Daemon_CP_1176_elements(43) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_1176_elements(40);
      outputPort_2_Daemon_CP_1176_elements(49)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(53);
      outputPort_2_Daemon_CP_1176_elements(50)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(54);
      outputPort_2_Daemon_CP_1176_elements(41) <= phi_mux_reqs(1);
      phi_stmt_883_phi_seq_1293 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_883_phi_seq_1293") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_1176_elements(36), 
          phi_sample_ack => outputPort_2_Daemon_CP_1176_elements(37), 
          phi_update_req => outputPort_2_Daemon_CP_1176_elements(38), 
          phi_update_ack => outputPort_2_Daemon_CP_1176_elements(39), 
          phi_mux_ack => outputPort_2_Daemon_CP_1176_elements(44), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_888_phi_seq_1337_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_1176_elements(63);
      outputPort_2_Daemon_CP_1176_elements(66)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(66);
      outputPort_2_Daemon_CP_1176_elements(67)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(68);
      outputPort_2_Daemon_CP_1176_elements(64) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_1176_elements(61);
      outputPort_2_Daemon_CP_1176_elements(70)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(74);
      outputPort_2_Daemon_CP_1176_elements(71)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(75);
      outputPort_2_Daemon_CP_1176_elements(62) <= phi_mux_reqs(1);
      phi_stmt_888_phi_seq_1337 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_888_phi_seq_1337") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_1176_elements(57), 
          phi_sample_ack => outputPort_2_Daemon_CP_1176_elements(58), 
          phi_update_req => outputPort_2_Daemon_CP_1176_elements(59), 
          phi_update_ack => outputPort_2_Daemon_CP_1176_elements(60), 
          phi_mux_ack => outputPort_2_Daemon_CP_1176_elements(65), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_893_phi_seq_1381_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_1176_elements(84);
      outputPort_2_Daemon_CP_1176_elements(87)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(87);
      outputPort_2_Daemon_CP_1176_elements(88)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(89);
      outputPort_2_Daemon_CP_1176_elements(85) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_1176_elements(82);
      outputPort_2_Daemon_CP_1176_elements(91)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(95);
      outputPort_2_Daemon_CP_1176_elements(92)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(96);
      outputPort_2_Daemon_CP_1176_elements(83) <= phi_mux_reqs(1);
      phi_stmt_893_phi_seq_1381 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_893_phi_seq_1381") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_1176_elements(78), 
          phi_sample_ack => outputPort_2_Daemon_CP_1176_elements(79), 
          phi_update_req => outputPort_2_Daemon_CP_1176_elements(80), 
          phi_update_ack => outputPort_2_Daemon_CP_1176_elements(81), 
          phi_mux_ack => outputPort_2_Daemon_CP_1176_elements(86), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_898_phi_seq_1425_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_1176_elements(105);
      outputPort_2_Daemon_CP_1176_elements(108)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(108);
      outputPort_2_Daemon_CP_1176_elements(109)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(110);
      outputPort_2_Daemon_CP_1176_elements(106) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_1176_elements(103);
      outputPort_2_Daemon_CP_1176_elements(112)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(116);
      outputPort_2_Daemon_CP_1176_elements(113)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(117);
      outputPort_2_Daemon_CP_1176_elements(104) <= phi_mux_reqs(1);
      phi_stmt_898_phi_seq_1425 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_898_phi_seq_1425") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_1176_elements(99), 
          phi_sample_ack => outputPort_2_Daemon_CP_1176_elements(100), 
          phi_update_req => outputPort_2_Daemon_CP_1176_elements(101), 
          phi_update_ack => outputPort_2_Daemon_CP_1176_elements(102), 
          phi_mux_ack => outputPort_2_Daemon_CP_1176_elements(107), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_903_phi_seq_1469_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_1176_elements(126);
      outputPort_2_Daemon_CP_1176_elements(129)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(129);
      outputPort_2_Daemon_CP_1176_elements(130)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(131);
      outputPort_2_Daemon_CP_1176_elements(127) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_1176_elements(124);
      outputPort_2_Daemon_CP_1176_elements(133)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(135);
      outputPort_2_Daemon_CP_1176_elements(134)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(136);
      outputPort_2_Daemon_CP_1176_elements(125) <= phi_mux_reqs(1);
      phi_stmt_903_phi_seq_1469 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_903_phi_seq_1469") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_1176_elements(120), 
          phi_sample_ack => outputPort_2_Daemon_CP_1176_elements(121), 
          phi_update_req => outputPort_2_Daemon_CP_1176_elements(122), 
          phi_update_ack => outputPort_2_Daemon_CP_1176_elements(123), 
          phi_mux_ack => outputPort_2_Daemon_CP_1176_elements(128), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_907_phi_seq_1513_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_2_Daemon_CP_1176_elements(143);
      outputPort_2_Daemon_CP_1176_elements(146)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(146);
      outputPort_2_Daemon_CP_1176_elements(147)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_2_Daemon_CP_1176_elements(148);
      outputPort_2_Daemon_CP_1176_elements(144) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_2_Daemon_CP_1176_elements(141);
      outputPort_2_Daemon_CP_1176_elements(150)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(152);
      outputPort_2_Daemon_CP_1176_elements(151)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_2_Daemon_CP_1176_elements(153);
      outputPort_2_Daemon_CP_1176_elements(142) <= phi_mux_reqs(1);
      phi_stmt_907_phi_seq_1513 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_907_phi_seq_1513") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_2_Daemon_CP_1176_elements(11), 
          phi_sample_ack => outputPort_2_Daemon_CP_1176_elements(139), 
          phi_update_req => outputPort_2_Daemon_CP_1176_elements(13), 
          phi_update_ack => outputPort_2_Daemon_CP_1176_elements(140), 
          phi_mux_ack => outputPort_2_Daemon_CP_1176_elements(145), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1201_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= outputPort_2_Daemon_CP_1176_elements(7);
        preds(1)  <= outputPort_2_Daemon_CP_1176_elements(8);
        entry_tmerge_1201 : transition_merge -- 
          generic map(name => " entry_tmerge_1201")
          port map (preds => preds, symbol_out => outputPort_2_Daemon_CP_1176_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u3_u1_1000_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1008_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1016_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1024_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1030_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1037_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1045_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1052_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1063_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1069_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1076_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1082_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_935_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_941_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_948_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_954_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_981_wire : std_logic_vector(0 downto 0);
    signal MUX_1034_wire : std_logic_vector(31 downto 0);
    signal MUX_1041_wire : std_logic_vector(31 downto 0);
    signal MUX_1049_wire : std_logic_vector(31 downto 0);
    signal MUX_1056_wire : std_logic_vector(31 downto 0);
    signal MUX_1066_wire : std_logic_vector(0 downto 0);
    signal MUX_1072_wire : std_logic_vector(0 downto 0);
    signal MUX_1079_wire : std_logic_vector(0 downto 0);
    signal MUX_1085_wire : std_logic_vector(0 downto 0);
    signal MUX_938_wire : std_logic_vector(0 downto 0);
    signal MUX_944_wire : std_logic_vector(0 downto 0);
    signal MUX_951_wire : std_logic_vector(0 downto 0);
    signal MUX_957_wire : std_logic_vector(0 downto 0);
    signal MUX_992_wire : std_logic_vector(7 downto 0);
    signal NOT_u1_u1_1005_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1013_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1021_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_997_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1073_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1086_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_945_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_958_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_974_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_977_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_978_wire : std_logic_vector(0 downto 0);
    signal OR_u32_u32_1042_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_1057_wire : std_logic_vector(31 downto 0);
    signal RPIPE_noblock_obuf_1_2_887_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_2_2_892_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_3_2_897_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_4_2_902_wire : std_logic_vector(32 downto 0);
    signal R_ZERO_33_885_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_890_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_895_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_900_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_3_905_wire_constant : std_logic_vector(2 downto 0);
    signal R_ZERO_3_909_wire_constant : std_logic_vector(2 downto 0);
    signal R_ZERO_8_881_wire_constant : std_logic_vector(7 downto 0);
    signal SUB_u8_u8_990_wire : std_logic_vector(7 downto 0);
    signal active_packet_903 : std_logic_vector(2 downto 0);
    signal data_to_out_1059 : std_logic_vector(31 downto 0);
    signal down_counter_879 : std_logic_vector(7 downto 0);
    signal konst_1007_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1015_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1023_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1029_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1033_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1036_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1040_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1044_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1048_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1051_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1055_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1062_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1065_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1068_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1071_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1075_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1078_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1081_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1084_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1094_wire_constant : std_logic_vector(0 downto 0);
    signal konst_914_wire_constant : std_logic_vector(32 downto 0);
    signal konst_919_wire_constant : std_logic_vector(32 downto 0);
    signal konst_924_wire_constant : std_logic_vector(32 downto 0);
    signal konst_929_wire_constant : std_logic_vector(32 downto 0);
    signal konst_934_wire_constant : std_logic_vector(2 downto 0);
    signal konst_937_wire_constant : std_logic_vector(0 downto 0);
    signal konst_940_wire_constant : std_logic_vector(2 downto 0);
    signal konst_943_wire_constant : std_logic_vector(0 downto 0);
    signal konst_947_wire_constant : std_logic_vector(2 downto 0);
    signal konst_950_wire_constant : std_logic_vector(0 downto 0);
    signal konst_953_wire_constant : std_logic_vector(2 downto 0);
    signal konst_956_wire_constant : std_logic_vector(0 downto 0);
    signal konst_980_wire_constant : std_logic_vector(7 downto 0);
    signal konst_986_wire_constant : std_logic_vector(7 downto 0);
    signal konst_989_wire_constant : std_logic_vector(7 downto 0);
    signal konst_999_wire_constant : std_logic_vector(2 downto 0);
    signal next_active_packet_970 : std_logic_vector(2 downto 0);
    signal next_active_packet_970_906_buffered : std_logic_vector(2 downto 0);
    signal next_down_counter_994 : std_logic_vector(7 downto 0);
    signal next_down_counter_994_882_buffered : std_logic_vector(7 downto 0);
    signal next_pkt_priority_970 : std_logic_vector(2 downto 0);
    signal next_pkt_priority_970_910_buffered : std_logic_vector(2 downto 0);
    signal p1_valid_916 : std_logic_vector(0 downto 0);
    signal p2_valid_921 : std_logic_vector(0 downto 0);
    signal p3_valid_926 : std_logic_vector(0 downto 0);
    signal p4_valid_931 : std_logic_vector(0 downto 0);
    signal pkt_1_e_word_883 : std_logic_vector(32 downto 0);
    signal pkt_2_e_word_888 : std_logic_vector(32 downto 0);
    signal pkt_3_e_word_893 : std_logic_vector(32 downto 0);
    signal pkt_4_e_word_898 : std_logic_vector(32 downto 0);
    signal pkt_priority_907 : std_logic_vector(2 downto 0);
    signal read_from_1_1002 : std_logic_vector(0 downto 0);
    signal read_from_2_1010 : std_logic_vector(0 downto 0);
    signal read_from_3_1018 : std_logic_vector(0 downto 0);
    signal read_from_4_1026 : std_logic_vector(0 downto 0);
    signal send_flag_1088 : std_logic_vector(0 downto 0);
    signal slice_1032_wire : std_logic_vector(31 downto 0);
    signal slice_1039_wire : std_logic_vector(31 downto 0);
    signal slice_1047_wire : std_logic_vector(31 downto 0);
    signal slice_1054_wire : std_logic_vector(31 downto 0);
    signal started_new_packet_983 : std_logic_vector(0 downto 0);
    signal valid_active_pkt_word_read_960 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_ZERO_33_885_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_890_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_895_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_900_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_3_905_wire_constant <= "000";
    R_ZERO_3_909_wire_constant <= "000";
    R_ZERO_8_881_wire_constant <= "00000000";
    konst_1007_wire_constant <= "010";
    konst_1015_wire_constant <= "011";
    konst_1023_wire_constant <= "100";
    konst_1029_wire_constant <= "001";
    konst_1033_wire_constant <= "00000000000000000000000000000000";
    konst_1036_wire_constant <= "010";
    konst_1040_wire_constant <= "00000000000000000000000000000000";
    konst_1044_wire_constant <= "011";
    konst_1048_wire_constant <= "00000000000000000000000000000000";
    konst_1051_wire_constant <= "100";
    konst_1055_wire_constant <= "00000000000000000000000000000000";
    konst_1062_wire_constant <= "001";
    konst_1065_wire_constant <= "0";
    konst_1068_wire_constant <= "010";
    konst_1071_wire_constant <= "0";
    konst_1075_wire_constant <= "011";
    konst_1078_wire_constant <= "0";
    konst_1081_wire_constant <= "100";
    konst_1084_wire_constant <= "0";
    konst_1094_wire_constant <= "1";
    konst_914_wire_constant <= "000000000000000000000000000100000";
    konst_919_wire_constant <= "000000000000000000000000000100000";
    konst_924_wire_constant <= "000000000000000000000000000100000";
    konst_929_wire_constant <= "000000000000000000000000000100000";
    konst_934_wire_constant <= "001";
    konst_937_wire_constant <= "0";
    konst_940_wire_constant <= "010";
    konst_943_wire_constant <= "0";
    konst_947_wire_constant <= "011";
    konst_950_wire_constant <= "0";
    konst_953_wire_constant <= "100";
    konst_956_wire_constant <= "0";
    konst_980_wire_constant <= "00000000";
    konst_986_wire_constant <= "00111111";
    konst_989_wire_constant <= "00000001";
    konst_999_wire_constant <= "001";
    phi_stmt_879: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_8_881_wire_constant & next_down_counter_994_882_buffered;
      req <= phi_stmt_879_req_0 & phi_stmt_879_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_879",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_879_ack_0,
          idata => idata,
          odata => down_counter_879,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_879
    phi_stmt_883: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_885_wire_constant & RPIPE_noblock_obuf_1_2_887_wire;
      req <= phi_stmt_883_req_0 & phi_stmt_883_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_883",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_883_ack_0,
          idata => idata,
          odata => pkt_1_e_word_883,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_883
    phi_stmt_888: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_890_wire_constant & RPIPE_noblock_obuf_2_2_892_wire;
      req <= phi_stmt_888_req_0 & phi_stmt_888_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_888",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_888_ack_0,
          idata => idata,
          odata => pkt_2_e_word_888,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_888
    phi_stmt_893: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_895_wire_constant & RPIPE_noblock_obuf_3_2_897_wire;
      req <= phi_stmt_893_req_0 & phi_stmt_893_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_893",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_893_ack_0,
          idata => idata,
          odata => pkt_3_e_word_893,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_893
    phi_stmt_898: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_900_wire_constant & RPIPE_noblock_obuf_4_2_902_wire;
      req <= phi_stmt_898_req_0 & phi_stmt_898_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_898",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_898_ack_0,
          idata => idata,
          odata => pkt_4_e_word_898,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_898
    phi_stmt_903: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_3_905_wire_constant & next_active_packet_970_906_buffered;
      req <= phi_stmt_903_req_0 & phi_stmt_903_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_903",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_903_ack_0,
          idata => idata,
          odata => active_packet_903,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_903
    phi_stmt_907: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_3_909_wire_constant & next_pkt_priority_970_910_buffered;
      req <= phi_stmt_907_req_0 & phi_stmt_907_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_907",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_907_ack_0,
          idata => idata,
          odata => pkt_priority_907,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_907
    -- flow-through select operator MUX_1034_inst
    MUX_1034_wire <= slice_1032_wire when (EQ_u3_u1_1030_wire(0) /=  '0') else konst_1033_wire_constant;
    -- flow-through select operator MUX_1041_inst
    MUX_1041_wire <= slice_1039_wire when (EQ_u3_u1_1037_wire(0) /=  '0') else konst_1040_wire_constant;
    -- flow-through select operator MUX_1049_inst
    MUX_1049_wire <= slice_1047_wire when (EQ_u3_u1_1045_wire(0) /=  '0') else konst_1048_wire_constant;
    -- flow-through select operator MUX_1056_inst
    MUX_1056_wire <= slice_1054_wire when (EQ_u3_u1_1052_wire(0) /=  '0') else konst_1055_wire_constant;
    -- flow-through select operator MUX_1066_inst
    MUX_1066_wire <= p1_valid_916 when (EQ_u3_u1_1063_wire(0) /=  '0') else konst_1065_wire_constant;
    -- flow-through select operator MUX_1072_inst
    MUX_1072_wire <= p2_valid_921 when (EQ_u3_u1_1069_wire(0) /=  '0') else konst_1071_wire_constant;
    -- flow-through select operator MUX_1079_inst
    MUX_1079_wire <= p3_valid_926 when (EQ_u3_u1_1076_wire(0) /=  '0') else konst_1078_wire_constant;
    -- flow-through select operator MUX_1085_inst
    MUX_1085_wire <= p4_valid_931 when (EQ_u3_u1_1082_wire(0) /=  '0') else konst_1084_wire_constant;
    -- flow-through select operator MUX_938_inst
    MUX_938_wire <= p1_valid_916 when (EQ_u3_u1_935_wire(0) /=  '0') else konst_937_wire_constant;
    -- flow-through select operator MUX_944_inst
    MUX_944_wire <= p2_valid_921 when (EQ_u3_u1_941_wire(0) /=  '0') else konst_943_wire_constant;
    -- flow-through select operator MUX_951_inst
    MUX_951_wire <= p3_valid_926 when (EQ_u3_u1_948_wire(0) /=  '0') else konst_950_wire_constant;
    -- flow-through select operator MUX_957_inst
    MUX_957_wire <= p4_valid_931 when (EQ_u3_u1_954_wire(0) /=  '0') else konst_956_wire_constant;
    -- flow-through select operator MUX_992_inst
    MUX_992_wire <= SUB_u8_u8_990_wire when (valid_active_pkt_word_read_960(0) /=  '0') else down_counter_879;
    -- flow-through select operator MUX_993_inst
    next_down_counter_994 <= konst_986_wire_constant when (started_new_packet_983(0) /=  '0') else MUX_992_wire;
    -- flow-through slice operator slice_1032_inst
    slice_1032_wire <= pkt_1_e_word_883(31 downto 0);
    -- flow-through slice operator slice_1039_inst
    slice_1039_wire <= pkt_2_e_word_888(31 downto 0);
    -- flow-through slice operator slice_1047_inst
    slice_1047_wire <= pkt_3_e_word_893(31 downto 0);
    -- flow-through slice operator slice_1054_inst
    slice_1054_wire <= pkt_4_e_word_898(31 downto 0);
    next_active_packet_970_906_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_active_packet_970_906_buf_req_0;
      next_active_packet_970_906_buf_ack_0<= wack(0);
      rreq(0) <= next_active_packet_970_906_buf_req_1;
      next_active_packet_970_906_buf_ack_1<= rack(0);
      next_active_packet_970_906_buf : InterlockBuffer generic map ( -- 
        name => "next_active_packet_970_906_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_active_packet_970,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_active_packet_970_906_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_down_counter_994_882_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_down_counter_994_882_buf_req_0;
      next_down_counter_994_882_buf_ack_0<= wack(0);
      rreq(0) <= next_down_counter_994_882_buf_req_1;
      next_down_counter_994_882_buf_ack_1<= rack(0);
      next_down_counter_994_882_buf : InterlockBuffer generic map ( -- 
        name => "next_down_counter_994_882_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_down_counter_994,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_down_counter_994_882_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_pkt_priority_970_910_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_pkt_priority_970_910_buf_req_0;
      next_pkt_priority_970_910_buf_ack_0<= wack(0);
      rreq(0) <= next_pkt_priority_970_910_buf_req_1;
      next_pkt_priority_970_910_buf_ack_1<= rack(0);
      next_pkt_priority_970_910_buf : InterlockBuffer generic map ( -- 
        name => "next_pkt_priority_970_910_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_pkt_priority_970,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_pkt_priority_970_910_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_877_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1094_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_877_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_877_branch_req_0,
          ack0 => do_while_stmt_877_branch_ack_0,
          ack1 => do_while_stmt_877_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator AND_u1_u1_982_inst
    process(OR_u1_u1_978_wire, EQ_u8_u1_981_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(OR_u1_u1_978_wire, EQ_u8_u1_981_wire, tmp_var);
      started_new_packet_983 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_915_inst
    process(pkt_1_e_word_883) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_1_e_word_883, konst_914_wire_constant, tmp_var);
      p1_valid_916 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_920_inst
    process(pkt_2_e_word_888) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_2_e_word_888, konst_919_wire_constant, tmp_var);
      p2_valid_921 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_925_inst
    process(pkt_3_e_word_893) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_3_e_word_893, konst_924_wire_constant, tmp_var);
      p3_valid_926 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_930_inst
    process(pkt_4_e_word_898) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_4_e_word_898, konst_929_wire_constant, tmp_var);
      p4_valid_931 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1000_inst
    process(next_active_packet_970) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_970, konst_999_wire_constant, tmp_var);
      EQ_u3_u1_1000_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1008_inst
    process(next_active_packet_970) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_970, konst_1007_wire_constant, tmp_var);
      EQ_u3_u1_1008_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1016_inst
    process(next_active_packet_970) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_970, konst_1015_wire_constant, tmp_var);
      EQ_u3_u1_1016_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1024_inst
    process(next_active_packet_970) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_970, konst_1023_wire_constant, tmp_var);
      EQ_u3_u1_1024_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1030_inst
    process(next_active_packet_970) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_970, konst_1029_wire_constant, tmp_var);
      EQ_u3_u1_1030_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1037_inst
    process(next_active_packet_970) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_970, konst_1036_wire_constant, tmp_var);
      EQ_u3_u1_1037_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1045_inst
    process(next_active_packet_970) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_970, konst_1044_wire_constant, tmp_var);
      EQ_u3_u1_1045_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1052_inst
    process(next_active_packet_970) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_970, konst_1051_wire_constant, tmp_var);
      EQ_u3_u1_1052_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1063_inst
    process(next_active_packet_970) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_970, konst_1062_wire_constant, tmp_var);
      EQ_u3_u1_1063_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1069_inst
    process(next_active_packet_970) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_970, konst_1068_wire_constant, tmp_var);
      EQ_u3_u1_1069_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1076_inst
    process(next_active_packet_970) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_970, konst_1075_wire_constant, tmp_var);
      EQ_u3_u1_1076_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1082_inst
    process(next_active_packet_970) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_970, konst_1081_wire_constant, tmp_var);
      EQ_u3_u1_1082_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_935_inst
    process(active_packet_903) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_903, konst_934_wire_constant, tmp_var);
      EQ_u3_u1_935_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_941_inst
    process(active_packet_903) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_903, konst_940_wire_constant, tmp_var);
      EQ_u3_u1_941_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_948_inst
    process(active_packet_903) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_903, konst_947_wire_constant, tmp_var);
      EQ_u3_u1_948_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_954_inst
    process(active_packet_903) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_903, konst_953_wire_constant, tmp_var);
      EQ_u3_u1_954_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_981_inst
    process(down_counter_879) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(down_counter_879, konst_980_wire_constant, tmp_var);
      EQ_u8_u1_981_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1005_inst
    process(p2_valid_921) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_921, tmp_var);
      NOT_u1_u1_1005_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1013_inst
    process(p3_valid_926) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_926, tmp_var);
      NOT_u1_u1_1013_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1021_inst
    process(p4_valid_931) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_931, tmp_var);
      NOT_u1_u1_1021_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_997_inst
    process(p1_valid_916) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_916, tmp_var);
      NOT_u1_u1_997_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1001_inst
    process(NOT_u1_u1_997_wire, EQ_u3_u1_1000_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_997_wire, EQ_u3_u1_1000_wire, tmp_var);
      read_from_1_1002 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1009_inst
    process(NOT_u1_u1_1005_wire, EQ_u3_u1_1008_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1005_wire, EQ_u3_u1_1008_wire, tmp_var);
      read_from_2_1010 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1017_inst
    process(NOT_u1_u1_1013_wire, EQ_u3_u1_1016_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1013_wire, EQ_u3_u1_1016_wire, tmp_var);
      read_from_3_1018 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1025_inst
    process(NOT_u1_u1_1021_wire, EQ_u3_u1_1024_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1021_wire, EQ_u3_u1_1024_wire, tmp_var);
      read_from_4_1026 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1073_inst
    process(MUX_1066_wire, MUX_1072_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1066_wire, MUX_1072_wire, tmp_var);
      OR_u1_u1_1073_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1086_inst
    process(MUX_1079_wire, MUX_1085_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1079_wire, MUX_1085_wire, tmp_var);
      OR_u1_u1_1086_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1087_inst
    process(OR_u1_u1_1073_wire, OR_u1_u1_1086_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1073_wire, OR_u1_u1_1086_wire, tmp_var);
      send_flag_1088 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_945_inst
    process(MUX_938_wire, MUX_944_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_938_wire, MUX_944_wire, tmp_var);
      OR_u1_u1_945_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_958_inst
    process(MUX_951_wire, MUX_957_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_951_wire, MUX_957_wire, tmp_var);
      OR_u1_u1_958_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_959_inst
    process(OR_u1_u1_945_wire, OR_u1_u1_958_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_945_wire, OR_u1_u1_958_wire, tmp_var);
      valid_active_pkt_word_read_960 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_974_inst
    process(p1_valid_916, p2_valid_921) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(p1_valid_916, p2_valid_921, tmp_var);
      OR_u1_u1_974_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_977_inst
    process(p3_valid_926, p4_valid_931) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(p3_valid_926, p4_valid_931, tmp_var);
      OR_u1_u1_977_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_978_inst
    process(OR_u1_u1_974_wire, OR_u1_u1_977_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_974_wire, OR_u1_u1_977_wire, tmp_var);
      OR_u1_u1_978_wire <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1042_inst
    process(MUX_1034_wire, MUX_1041_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1034_wire, MUX_1041_wire, tmp_var);
      OR_u32_u32_1042_wire <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1057_inst
    process(MUX_1049_wire, MUX_1056_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1049_wire, MUX_1056_wire, tmp_var);
      OR_u32_u32_1057_wire <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1058_inst
    process(OR_u32_u32_1042_wire, OR_u32_u32_1057_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u32_u32_1042_wire, OR_u32_u32_1057_wire, tmp_var);
      data_to_out_1059 <= tmp_var; --
    end process;
    -- binary operator SUB_u8_u8_990_inst
    process(down_counter_879) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSub_proc(down_counter_879, konst_989_wire_constant, tmp_var);
      SUB_u8_u8_990_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_noblock_obuf_1_2_887_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_1_2_887_inst_req_0;
      RPIPE_noblock_obuf_1_2_887_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_1_2_887_inst_req_1;
      RPIPE_noblock_obuf_1_2_887_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_1_1002(0);
      RPIPE_noblock_obuf_1_2_887_wire <= data_out(32 downto 0);
      noblock_obuf_1_2_read_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_2_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_2_read_0: InputPortRevised -- 
        generic map ( name => "noblock_obuf_1_2_read_0", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_1_2_pipe_read_req(0),
          oack => noblock_obuf_1_2_pipe_read_ack(0),
          odata => noblock_obuf_1_2_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_noblock_obuf_2_2_892_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_2_2_892_inst_req_0;
      RPIPE_noblock_obuf_2_2_892_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_2_2_892_inst_req_1;
      RPIPE_noblock_obuf_2_2_892_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_2_1010(0);
      RPIPE_noblock_obuf_2_2_892_wire <= data_out(32 downto 0);
      noblock_obuf_2_2_read_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_2_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_2_read_1: InputPortRevised -- 
        generic map ( name => "noblock_obuf_2_2_read_1", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_2_2_pipe_read_req(0),
          oack => noblock_obuf_2_2_pipe_read_ack(0),
          odata => noblock_obuf_2_2_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_noblock_obuf_3_2_897_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_3_2_897_inst_req_0;
      RPIPE_noblock_obuf_3_2_897_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_3_2_897_inst_req_1;
      RPIPE_noblock_obuf_3_2_897_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_3_1018(0);
      RPIPE_noblock_obuf_3_2_897_wire <= data_out(32 downto 0);
      noblock_obuf_3_2_read_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_2_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_2_read_2: InputPortRevised -- 
        generic map ( name => "noblock_obuf_3_2_read_2", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_3_2_pipe_read_req(0),
          oack => noblock_obuf_3_2_pipe_read_ack(0),
          odata => noblock_obuf_3_2_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_noblock_obuf_4_2_902_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_4_2_902_inst_req_0;
      RPIPE_noblock_obuf_4_2_902_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_4_2_902_inst_req_1;
      RPIPE_noblock_obuf_4_2_902_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_4_1026(0);
      RPIPE_noblock_obuf_4_2_902_wire <= data_out(32 downto 0);
      noblock_obuf_4_2_read_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_2_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_2_read_3: InputPortRevised -- 
        generic map ( name => "noblock_obuf_4_2_read_3", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_4_2_pipe_read_req(0),
          oack => noblock_obuf_4_2_pipe_read_ack(0),
          odata => noblock_obuf_4_2_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_out_data_2_1090_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_out_data_2_1090_inst_req_0;
      WPIPE_out_data_2_1090_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_out_data_2_1090_inst_req_1;
      WPIPE_out_data_2_1090_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_flag_1088(0);
      data_in <= data_to_out_1059;
      out_data_2_write_0_gI: SplitGuardInterface generic map(name => "out_data_2_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      out_data_2_write_0: OutputPortRevised -- 
        generic map ( name => "out_data_2", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => out_data_2_pipe_write_req(0),
          oack => out_data_2_pipe_write_ack(0),
          odata => out_data_2_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    volatile_operator_prioritySelect_2575: prioritySelect_Volatile port map(down_counter => down_counter_879, active_packet => active_packet_903, pkt_priority => pkt_priority_907, p1_valid => p1_valid_916, p2_valid => p2_valid_921, p3_valid => p3_valid_926, p4_valid => p4_valid_931, next_active_packet => next_active_packet_970, next_pkt_priority => next_pkt_priority_970); 
    -- 
  end Block; -- data_path
  -- 
end outputPort_2_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity outputPort_3_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    noblock_obuf_1_3_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_3_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_3_3_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_3_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_4_3_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_3_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_2_3_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_3_pipe_read_data : in   std_logic_vector(32 downto 0);
    out_data_3_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_3_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity outputPort_3_Daemon;
architecture outputPort_3_Daemon_arch of outputPort_3_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal outputPort_3_Daemon_CP_1538_start: Boolean;
  signal outputPort_3_Daemon_CP_1538_symbol: Boolean;
  -- volatile/operator module components. 
  component prioritySelect_Volatile is -- 
    port ( -- 
      down_counter : in  std_logic_vector(7 downto 0);
      active_packet : in  std_logic_vector(2 downto 0);
      pkt_priority : in  std_logic_vector(2 downto 0);
      p1_valid : in  std_logic_vector(0 downto 0);
      p2_valid : in  std_logic_vector(0 downto 0);
      p3_valid : in  std_logic_vector(0 downto 0);
      p4_valid : in  std_logic_vector(0 downto 0);
      next_active_packet : out  std_logic_vector(2 downto 0);
      next_pkt_priority : out  std_logic_vector(2 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal RPIPE_noblock_obuf_1_3_1109_inst_ack_1 : boolean;
  signal phi_stmt_1110_req_1 : boolean;
  signal next_down_counter_1216_1104_buf_ack_1 : boolean;
  signal phi_stmt_1110_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_3_1109_inst_ack_0 : boolean;
  signal phi_stmt_1110_req_0 : boolean;
  signal do_while_stmt_1099_branch_req_0 : boolean;
  signal phi_stmt_1105_ack_0 : boolean;
  signal next_down_counter_1216_1104_buf_req_1 : boolean;
  signal RPIPE_noblock_obuf_3_3_1119_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_3_3_1119_inst_ack_1 : boolean;
  signal next_active_packet_1192_1128_buf_req_0 : boolean;
  signal next_active_packet_1192_1128_buf_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_3_1109_inst_req_0 : boolean;
  signal next_down_counter_1216_1104_buf_req_0 : boolean;
  signal next_down_counter_1216_1104_buf_ack_0 : boolean;
  signal RPIPE_noblock_obuf_1_3_1109_inst_req_1 : boolean;
  signal phi_stmt_1125_req_1 : boolean;
  signal RPIPE_noblock_obuf_4_3_1124_inst_ack_1 : boolean;
  signal RPIPE_noblock_obuf_4_3_1124_inst_req_1 : boolean;
  signal phi_stmt_1120_ack_0 : boolean;
  signal phi_stmt_1120_req_0 : boolean;
  signal phi_stmt_1125_req_0 : boolean;
  signal phi_stmt_1101_ack_0 : boolean;
  signal RPIPE_noblock_obuf_4_3_1124_inst_ack_0 : boolean;
  signal phi_stmt_1120_req_1 : boolean;
  signal RPIPE_noblock_obuf_4_3_1124_inst_req_0 : boolean;
  signal phi_stmt_1101_req_0 : boolean;
  signal phi_stmt_1101_req_1 : boolean;
  signal RPIPE_noblock_obuf_2_3_1114_inst_ack_0 : boolean;
  signal phi_stmt_1129_req_1 : boolean;
  signal RPIPE_noblock_obuf_2_3_1114_inst_req_0 : boolean;
  signal phi_stmt_1129_req_0 : boolean;
  signal RPIPE_noblock_obuf_3_3_1119_inst_ack_0 : boolean;
  signal phi_stmt_1115_ack_0 : boolean;
  signal RPIPE_noblock_obuf_3_3_1119_inst_req_0 : boolean;
  signal next_active_packet_1192_1128_buf_ack_1 : boolean;
  signal phi_stmt_1115_req_0 : boolean;
  signal phi_stmt_1115_req_1 : boolean;
  signal phi_stmt_1129_ack_0 : boolean;
  signal phi_stmt_1105_req_0 : boolean;
  signal next_active_packet_1192_1128_buf_req_1 : boolean;
  signal phi_stmt_1105_req_1 : boolean;
  signal RPIPE_noblock_obuf_2_3_1114_inst_ack_1 : boolean;
  signal phi_stmt_1125_ack_0 : boolean;
  signal RPIPE_noblock_obuf_2_3_1114_inst_req_1 : boolean;
  signal next_pkt_priority_1192_1132_buf_req_0 : boolean;
  signal next_pkt_priority_1192_1132_buf_ack_0 : boolean;
  signal next_pkt_priority_1192_1132_buf_req_1 : boolean;
  signal next_pkt_priority_1192_1132_buf_ack_1 : boolean;
  signal WPIPE_out_data_3_1312_inst_req_0 : boolean;
  signal WPIPE_out_data_3_1312_inst_ack_0 : boolean;
  signal WPIPE_out_data_3_1312_inst_req_1 : boolean;
  signal WPIPE_out_data_3_1312_inst_ack_1 : boolean;
  signal do_while_stmt_1099_branch_ack_0 : boolean;
  signal do_while_stmt_1099_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "outputPort_3_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  outputPort_3_Daemon_CP_1538_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "outputPort_3_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_3_Daemon_CP_1538_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= outputPort_3_Daemon_CP_1538_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_3_Daemon_CP_1538_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  outputPort_3_Daemon_CP_1538: Block -- control-path 
    signal outputPort_3_Daemon_CP_1538_elements: BooleanArray(161 downto 0);
    -- 
  begin -- 
    outputPort_3_Daemon_CP_1538_elements(0) <= outputPort_3_Daemon_CP_1538_start;
    outputPort_3_Daemon_CP_1538_symbol <= outputPort_3_Daemon_CP_1538_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1098/do_while_stmt_1099__entry__
      -- CP-element group 0: 	 branch_block_stmt_1098/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1098/branch_block_stmt_1098__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	161 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1098/do_while_stmt_1099__exit__
      -- CP-element group 1: 	 branch_block_stmt_1098/branch_block_stmt_1098__exit__
      -- CP-element group 1: 	 branch_block_stmt_1098/$exit
      -- CP-element group 1: 	 $exit
      -- 
    outputPort_3_Daemon_CP_1538_elements(1) <= outputPort_3_Daemon_CP_1538_elements(161);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099__entry__
      -- CP-element group 2: 	 branch_block_stmt_1098/do_while_stmt_1099/$entry
      -- 
    outputPort_3_Daemon_CP_1538_elements(2) <= outputPort_3_Daemon_CP_1538_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	161 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099__exit__
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1098/do_while_stmt_1099/loop_back
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	159 
    -- CP-element group 5: 	160 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1098/do_while_stmt_1099/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1098/do_while_stmt_1099/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1098/do_while_stmt_1099/loop_taken/$entry
      -- 
    outputPort_3_Daemon_CP_1538_elements(5) <= outputPort_3_Daemon_CP_1538_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	158 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1098/do_while_stmt_1099/loop_body_done
      -- 
    outputPort_3_Daemon_CP_1538_elements(6) <= outputPort_3_Daemon_CP_1538_elements(158);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	122 
    -- CP-element group 7: 	61 
    -- CP-element group 7: 	103 
    -- CP-element group 7: 	82 
    -- CP-element group 7: 	141 
    -- CP-element group 7: 	21 
    -- CP-element group 7: 	40 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/back_edge_to_loop_body
      -- 
    outputPort_3_Daemon_CP_1538_elements(7) <= outputPort_3_Daemon_CP_1538_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	63 
    -- CP-element group 8: 	105 
    -- CP-element group 8: 	124 
    -- CP-element group 8: 	84 
    -- CP-element group 8: 	143 
    -- CP-element group 8: 	23 
    -- CP-element group 8: 	42 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/first_time_through_loop_body
      -- 
    outputPort_3_Daemon_CP_1538_elements(8) <= outputPort_3_Daemon_CP_1538_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	118 
    -- CP-element group 9: 	119 
    -- CP-element group 9: 	157 
    -- CP-element group 9: 	76 
    -- CP-element group 9: 	135 
    -- CP-element group 9: 	136 
    -- CP-element group 9: 	97 
    -- CP-element group 9: 	55 
    -- CP-element group 9: 	56 
    -- CP-element group 9: 	98 
    -- CP-element group 9: 	77 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	34 
    -- CP-element group 9: 	35 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/loop_body_start
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	157 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/condition_evaluated
      -- 
    condition_evaluated_1562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(10), ack => do_while_stmt_1099_branch_req_0); -- 
    outputPort_3_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(157) & outputPort_3_Daemon_CP_1538_elements(14);
      gj_outputPort_3_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	118 
    -- CP-element group 11: 	76 
    -- CP-element group 11: 	135 
    -- CP-element group 11: 	97 
    -- CP-element group 11: 	55 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	34 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	78 
    -- CP-element group 11: 	57 
    -- CP-element group 11: 	99 
    -- CP-element group 11: 	137 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	36 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1125_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/aggregated_phi_sample_req
      -- 
    outputPort_3_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(118) & outputPort_3_Daemon_CP_1538_elements(76) & outputPort_3_Daemon_CP_1538_elements(135) & outputPort_3_Daemon_CP_1538_elements(97) & outputPort_3_Daemon_CP_1538_elements(55) & outputPort_3_Daemon_CP_1538_elements(15) & outputPort_3_Daemon_CP_1538_elements(34) & outputPort_3_Daemon_CP_1538_elements(14);
      gj_outputPort_3_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	120 
    -- CP-element group 12: 	100 
    -- CP-element group 12: 	79 
    -- CP-element group 12: 	58 
    -- CP-element group 12: 	138 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	37 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	158 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	118 
    -- CP-element group 12: 	76 
    -- CP-element group 12: 	135 
    -- CP-element group 12: 	97 
    -- CP-element group 12: 	55 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	34 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1101_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1105_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1115_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1110_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1120_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1125_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1129_sample_completed_
      -- 
    outputPort_3_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(120) & outputPort_3_Daemon_CP_1538_elements(100) & outputPort_3_Daemon_CP_1538_elements(79) & outputPort_3_Daemon_CP_1538_elements(58) & outputPort_3_Daemon_CP_1538_elements(138) & outputPort_3_Daemon_CP_1538_elements(18) & outputPort_3_Daemon_CP_1538_elements(37);
      gj_outputPort_3_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	119 
    -- CP-element group 13: 	136 
    -- CP-element group 13: 	56 
    -- CP-element group 13: 	98 
    -- CP-element group 13: 	77 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	35 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	101 
    -- CP-element group 13: 	59 
    -- CP-element group 13: 	80 
    -- CP-element group 13: 	139 
    -- CP-element group 13: 	19 
    -- CP-element group 13: 	38 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1125_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/aggregated_phi_update_req
      -- 
    outputPort_3_Daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(119) & outputPort_3_Daemon_CP_1538_elements(136) & outputPort_3_Daemon_CP_1538_elements(56) & outputPort_3_Daemon_CP_1538_elements(98) & outputPort_3_Daemon_CP_1538_elements(77) & outputPort_3_Daemon_CP_1538_elements(16) & outputPort_3_Daemon_CP_1538_elements(35);
      gj_outputPort_3_Daemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	121 
    -- CP-element group 14: 	102 
    -- CP-element group 14: 	60 
    -- CP-element group 14: 	81 
    -- CP-element group 14: 	140 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	39 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/aggregated_phi_update_ack
      -- 
    outputPort_3_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(121) & outputPort_3_Daemon_CP_1538_elements(102) & outputPort_3_Daemon_CP_1538_elements(60) & outputPort_3_Daemon_CP_1538_elements(81) & outputPort_3_Daemon_CP_1538_elements(140) & outputPort_3_Daemon_CP_1538_elements(20) & outputPort_3_Daemon_CP_1538_elements(39);
      gj_outputPort_3_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1101_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	155 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1101_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(155);
      gj_outputPort_3_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1101_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(17) <= outputPort_3_Daemon_CP_1538_elements(11);
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1101_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1101_update_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(19) <= outputPort_3_Daemon_CP_1538_elements(13);
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	154 
    -- CP-element group 20: 	14 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1101_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1101_update_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1101_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(21) <= outputPort_3_Daemon_CP_1538_elements(7);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1101_loopback_sample_req_ps
      -- CP-element group 22: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1101_loopback_sample_req
      -- 
    phi_stmt_1101_loopback_sample_req_1577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1101_loopback_sample_req_1577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(22), ack => phi_stmt_1101_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1101_entry_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(23) <= outputPort_3_Daemon_CP_1538_elements(8);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1101_entry_sample_req_ps
      -- CP-element group 24: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1101_entry_sample_req
      -- 
    phi_stmt_1101_entry_sample_req_1580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1101_entry_sample_req_1580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(24), ack => phi_stmt_1101_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1101_phi_mux_ack_ps
      -- CP-element group 25: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1101_phi_mux_ack
      -- 
    phi_stmt_1101_phi_mux_ack_1583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1101_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_8_1103_sample_start__ps
      -- CP-element group 26: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_8_1103_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_8_1103_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_8_1103_sample_start_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_8_1103_update_start_
      -- CP-element group 27: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_8_1103_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_8_1103_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(28) <= outputPort_3_Daemon_CP_1538_elements(29);
    -- CP-element group 29:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	28 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_8_1103_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(29) is a control-delay.
    cp_element_29_delay: control_delay_element  generic map(name => " 29_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_1538_elements(27), ack => outputPort_3_Daemon_CP_1538_elements(29), clk => clk, reset =>reset);
    -- CP-element group 30:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_down_counter_1104_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_down_counter_1104_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_down_counter_1104_Sample/req
      -- CP-element group 30: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_down_counter_1104_sample_start__ps
      -- 
    req_1604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(30), ack => next_down_counter_1216_1104_buf_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_down_counter_1104_Update/req
      -- CP-element group 31: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_down_counter_1104_update_start_
      -- CP-element group 31: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_down_counter_1104_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_down_counter_1104_update_start__ps
      -- 
    req_1609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(31), ack => next_down_counter_1216_1104_buf_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_down_counter_1104_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_down_counter_1104_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_down_counter_1104_Sample/ack
      -- CP-element group 32: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_down_counter_1104_sample_completed__ps
      -- 
    ack_1605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_1216_1104_buf_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(32)); -- 
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_down_counter_1104_Update/ack
      -- CP-element group 33: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_down_counter_1104_update_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_down_counter_1104_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_down_counter_1104_update_completed_
      -- 
    ack_1610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_1216_1104_buf_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(33)); -- 
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	9 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	12 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	11 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1105_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	155 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	13 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1105_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(155);
      gj_outputPort_3_Daemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	11 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1105_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(36) <= outputPort_3_Daemon_CP_1538_elements(11);
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	12 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1105_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1105_update_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(38) <= outputPort_3_Daemon_CP_1538_elements(13);
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	154 
    -- CP-element group 39: 	14 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1105_update_completed__ps
      -- CP-element group 39: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1105_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	7 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1105_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(40) <= outputPort_3_Daemon_CP_1538_elements(7);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1105_loopback_sample_req_ps
      -- CP-element group 41: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1105_loopback_sample_req
      -- 
    phi_stmt_1105_loopback_sample_req_1621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1105_loopback_sample_req_1621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(41), ack => phi_stmt_1105_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	8 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1105_entry_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(42) <= outputPort_3_Daemon_CP_1538_elements(8);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1105_entry_sample_req_ps
      -- CP-element group 43: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1105_entry_sample_req
      -- 
    phi_stmt_1105_entry_sample_req_1624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1105_entry_sample_req_1624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(43), ack => phi_stmt_1105_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1105_phi_mux_ack
      -- CP-element group 44: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1105_phi_mux_ack_ps
      -- 
    phi_stmt_1105_phi_mux_ack_1627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1105_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1107_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1107_sample_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1107_sample_start__ps
      -- CP-element group 45: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1107_sample_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1107_update_start__ps
      -- CP-element group 46: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1107_update_start_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1107_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(47) <= outputPort_3_Daemon_CP_1538_elements(48);
    -- CP-element group 48:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	47 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1107_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(48) is a control-delay.
    cp_element_48_delay: control_delay_element  generic map(name => " 48_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_1538_elements(46), ack => outputPort_3_Daemon_CP_1538_elements(48), clk => clk, reset =>reset);
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_1_3_1109_sample_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_1_3_1109_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	54 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_1_3_1109_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_1_3_1109_Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_1_3_1109_Sample/$entry
      -- 
    rr_1648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(51), ack => RPIPE_noblock_obuf_1_3_1109_inst_req_0); -- 
    outputPort_3_Daemon_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(49) & outputPort_3_Daemon_CP_1538_elements(54);
      gj_outputPort_3_Daemon_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	53 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_1_3_1109_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_1_3_1109_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_1_3_1109_Update/cr
      -- 
    cr_1653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(52), ack => RPIPE_noblock_obuf_1_3_1109_inst_req_1); -- 
    outputPort_3_Daemon_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(53) & outputPort_3_Daemon_CP_1538_elements(50);
      gj_outputPort_3_Daemon_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	52 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_1_3_1109_sample_completed__ps
      -- CP-element group 53: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_1_3_1109_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_1_3_1109_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_1_3_1109_Sample/$exit
      -- 
    ra_1649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_3_1109_inst_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(53)); -- 
    -- CP-element group 54:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	51 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_1_3_1109_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_1_3_1109_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_1_3_1109_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_1_3_1109_update_completed__ps
      -- 
    ca_1654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_3_1109_inst_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(54)); -- 
    -- CP-element group 55:  join  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	9 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	12 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	11 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1110_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	9 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	155 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	13 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1110_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(155);
      gj_outputPort_3_Daemon_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	11 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1110_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(57) <= outputPort_3_Daemon_CP_1538_elements(11);
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	12 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1110_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	13 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1110_update_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(59) <= outputPort_3_Daemon_CP_1538_elements(13);
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	154 
    -- CP-element group 60: 	14 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1110_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1110_update_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	7 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1110_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(61) <= outputPort_3_Daemon_CP_1538_elements(7);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1110_loopback_sample_req
      -- CP-element group 62: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1110_loopback_sample_req_ps
      -- 
    phi_stmt_1110_loopback_sample_req_1665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1110_loopback_sample_req_1665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(62), ack => phi_stmt_1110_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	8 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1110_entry_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(63) <= outputPort_3_Daemon_CP_1538_elements(8);
    -- CP-element group 64:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1110_entry_sample_req_ps
      -- CP-element group 64: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1110_entry_sample_req
      -- 
    phi_stmt_1110_entry_sample_req_1668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1110_entry_sample_req_1668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(64), ack => phi_stmt_1110_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1110_phi_mux_ack
      -- CP-element group 65: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1110_phi_mux_ack_ps
      -- 
    phi_stmt_1110_phi_mux_ack_1671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1110_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(65)); -- 
    -- CP-element group 66:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1112_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1112_sample_completed__ps
      -- CP-element group 66: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1112_sample_start__ps
      -- CP-element group 66: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1112_sample_start_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1112_update_start__ps
      -- CP-element group 67: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1112_update_start_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1112_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(68) <= outputPort_3_Daemon_CP_1538_elements(69);
    -- CP-element group 69:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	68 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1112_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(69) is a control-delay.
    cp_element_69_delay: control_delay_element  generic map(name => " 69_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_1538_elements(67), ack => outputPort_3_Daemon_CP_1538_elements(69), clk => clk, reset =>reset);
    -- CP-element group 70:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_2_3_1114_sample_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(70) is bound as output of CP function.
    -- CP-element group 71:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_2_3_1114_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: marked-predecessors 
    -- CP-element group 72: 	75 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_2_3_1114_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_2_3_1114_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_2_3_1114_Sample/rr
      -- 
    rr_1692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(72), ack => RPIPE_noblock_obuf_2_3_1114_inst_req_0); -- 
    outputPort_3_Daemon_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(70) & outputPort_3_Daemon_CP_1538_elements(75);
      gj_outputPort_3_Daemon_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	74 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_2_3_1114_update_start_
      -- CP-element group 73: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_2_3_1114_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_2_3_1114_Update/cr
      -- 
    cr_1697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(73), ack => RPIPE_noblock_obuf_2_3_1114_inst_req_1); -- 
    outputPort_3_Daemon_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(74) & outputPort_3_Daemon_CP_1538_elements(71);
      gj_outputPort_3_Daemon_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	73 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_2_3_1114_sample_completed__ps
      -- CP-element group 74: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_2_3_1114_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_2_3_1114_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_2_3_1114_Sample/ra
      -- 
    ra_1693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_3_1114_inst_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(74)); -- 
    -- CP-element group 75:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	72 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_2_3_1114_update_completed__ps
      -- CP-element group 75: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_2_3_1114_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_2_3_1114_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_2_3_1114_Update/ca
      -- 
    ca_1698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_3_1114_inst_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(75)); -- 
    -- CP-element group 76:  join  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	9 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	12 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	11 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1115_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	9 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	155 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	13 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1115_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(155);
      gj_outputPort_3_Daemon_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	11 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1115_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(78) <= outputPort_3_Daemon_CP_1538_elements(11);
    -- CP-element group 79:  join  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	12 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1115_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	13 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1115_update_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(80) <= outputPort_3_Daemon_CP_1538_elements(13);
    -- CP-element group 81:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	154 
    -- CP-element group 81: 	14 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1115_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1115_update_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	7 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1115_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(82) <= outputPort_3_Daemon_CP_1538_elements(7);
    -- CP-element group 83:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1115_loopback_sample_req_ps
      -- CP-element group 83: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1115_loopback_sample_req
      -- 
    phi_stmt_1115_loopback_sample_req_1709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1115_loopback_sample_req_1709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(83), ack => phi_stmt_1115_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(83) is bound as output of CP function.
    -- CP-element group 84:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	8 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1115_entry_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(84) <= outputPort_3_Daemon_CP_1538_elements(8);
    -- CP-element group 85:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1115_entry_sample_req_ps
      -- CP-element group 85: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1115_entry_sample_req
      -- 
    phi_stmt_1115_entry_sample_req_1712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1115_entry_sample_req_1712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(85), ack => phi_stmt_1115_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1115_phi_mux_ack_ps
      -- CP-element group 86: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1115_phi_mux_ack
      -- 
    phi_stmt_1115_phi_mux_ack_1715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1115_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(86)); -- 
    -- CP-element group 87:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1117_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1117_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1117_sample_completed__ps
      -- CP-element group 87: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1117_sample_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1117_update_start__ps
      -- CP-element group 88: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1117_update_start_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	90 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1117_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(89) <= outputPort_3_Daemon_CP_1538_elements(90);
    -- CP-element group 90:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	89 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1117_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(90) is a control-delay.
    cp_element_90_delay: control_delay_element  generic map(name => " 90_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_1538_elements(88), ack => outputPort_3_Daemon_CP_1538_elements(90), clk => clk, reset =>reset);
    -- CP-element group 91:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_3_3_1119_sample_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(91) is bound as output of CP function.
    -- CP-element group 92:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_3_3_1119_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(92) is bound as output of CP function.
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	96 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_3_3_1119_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_3_3_1119_Sample/rr
      -- CP-element group 93: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_3_3_1119_Sample/$entry
      -- 
    rr_1736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(93), ack => RPIPE_noblock_obuf_3_3_1119_inst_req_0); -- 
    outputPort_3_Daemon_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(91) & outputPort_3_Daemon_CP_1538_elements(96);
      gj_outputPort_3_Daemon_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	95 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_3_3_1119_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_3_3_1119_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_3_3_1119_Update/$entry
      -- 
    cr_1741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(94), ack => RPIPE_noblock_obuf_3_3_1119_inst_req_1); -- 
    outputPort_3_Daemon_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(92) & outputPort_3_Daemon_CP_1538_elements(95);
      gj_outputPort_3_Daemon_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	94 
    -- CP-element group 95:  members (4) 
      -- CP-element group 95: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_3_3_1119_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_3_3_1119_sample_completed__ps
      -- CP-element group 95: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_3_3_1119_Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_3_3_1119_Sample/$exit
      -- 
    ra_1737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_3_1119_inst_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(95)); -- 
    -- CP-element group 96:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	93 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_3_3_1119_Update/ca
      -- CP-element group 96: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_3_3_1119_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_3_3_1119_update_completed__ps
      -- CP-element group 96: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_3_3_1119_Update/$exit
      -- 
    ca_1742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_3_1119_inst_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(96)); -- 
    -- CP-element group 97:  join  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	9 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	12 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	11 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1120_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	9 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	155 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	13 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1120_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_3_Daemon_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(155);
      gj_outputPort_3_Daemon_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	11 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1120_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(99) <= outputPort_3_Daemon_CP_1538_elements(11);
    -- CP-element group 100:  join  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	12 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1120_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(100) is bound as output of CP function.
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	13 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1120_update_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(101) <= outputPort_3_Daemon_CP_1538_elements(13);
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	154 
    -- CP-element group 102: 	14 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1120_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1120_update_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(102) is bound as output of CP function.
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	7 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1120_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(103) <= outputPort_3_Daemon_CP_1538_elements(7);
    -- CP-element group 104:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1120_loopback_sample_req_ps
      -- CP-element group 104: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1120_loopback_sample_req
      -- 
    phi_stmt_1120_loopback_sample_req_1753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1120_loopback_sample_req_1753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(104), ack => phi_stmt_1120_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(104) is bound as output of CP function.
    -- CP-element group 105:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	8 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1120_entry_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(105) <= outputPort_3_Daemon_CP_1538_elements(8);
    -- CP-element group 106:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1120_entry_sample_req_ps
      -- CP-element group 106: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1120_entry_sample_req
      -- 
    phi_stmt_1120_entry_sample_req_1756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1120_entry_sample_req_1756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(106), ack => phi_stmt_1120_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1120_phi_mux_ack_ps
      -- CP-element group 107: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1120_phi_mux_ack
      -- 
    phi_stmt_1120_phi_mux_ack_1759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1120_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(107)); -- 
    -- CP-element group 108:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1122_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1122_sample_completed__ps
      -- CP-element group 108: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1122_sample_start__ps
      -- CP-element group 108: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1122_sample_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(108) is bound as output of CP function.
    -- CP-element group 109:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1122_update_start_
      -- CP-element group 109: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1122_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	111 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1122_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(110) <= outputPort_3_Daemon_CP_1538_elements(111);
    -- CP-element group 111:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	110 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_33_1122_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(111) is a control-delay.
    cp_element_111_delay: control_delay_element  generic map(name => " 111_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_1538_elements(109), ack => outputPort_3_Daemon_CP_1538_elements(111), clk => clk, reset =>reset);
    -- CP-element group 112:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_4_3_1124_sample_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(112) is bound as output of CP function.
    -- CP-element group 113:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_4_3_1124_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(113) is bound as output of CP function.
    -- CP-element group 114:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: marked-predecessors 
    -- CP-element group 114: 	117 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_4_3_1124_Sample/rr
      -- CP-element group 114: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_4_3_1124_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_4_3_1124_sample_start_
      -- 
    rr_1780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(114), ack => RPIPE_noblock_obuf_4_3_1124_inst_req_0); -- 
    outputPort_3_Daemon_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(112) & outputPort_3_Daemon_CP_1538_elements(117);
      gj_outputPort_3_Daemon_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	116 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_4_3_1124_Update/cr
      -- CP-element group 115: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_4_3_1124_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_4_3_1124_update_start_
      -- 
    cr_1785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(115), ack => RPIPE_noblock_obuf_4_3_1124_inst_req_1); -- 
    outputPort_3_Daemon_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(116) & outputPort_3_Daemon_CP_1538_elements(113);
      gj_outputPort_3_Daemon_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	115 
    -- CP-element group 116:  members (4) 
      -- CP-element group 116: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_4_3_1124_sample_completed__ps
      -- CP-element group 116: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_4_3_1124_Sample/ra
      -- CP-element group 116: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_4_3_1124_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_4_3_1124_sample_completed_
      -- 
    ra_1781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_3_1124_inst_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(116)); -- 
    -- CP-element group 117:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: marked-successors 
    -- CP-element group 117: 	114 
    -- CP-element group 117:  members (4) 
      -- CP-element group 117: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_4_3_1124_Update/ca
      -- CP-element group 117: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_4_3_1124_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_4_3_1124_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/RPIPE_noblock_obuf_4_3_1124_update_completed__ps
      -- 
    ca_1786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_3_1124_inst_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(117)); -- 
    -- CP-element group 118:  join  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	9 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	12 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	11 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1125_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  join  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	9 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	155 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	13 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1125_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(155);
      gj_outputPort_3_Daemon_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  join  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	12 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1125_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(120) is bound as output of CP function.
    -- CP-element group 121:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	154 
    -- CP-element group 121: 	14 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1125_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1125_update_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(121) is bound as output of CP function.
    -- CP-element group 122:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	7 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1125_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(122) <= outputPort_3_Daemon_CP_1538_elements(7);
    -- CP-element group 123:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1125_loopback_sample_req_ps
      -- CP-element group 123: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1125_loopback_sample_req
      -- 
    phi_stmt_1125_loopback_sample_req_1797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1125_loopback_sample_req_1797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(123), ack => phi_stmt_1125_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(123) is bound as output of CP function.
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	8 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1125_entry_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(124) <= outputPort_3_Daemon_CP_1538_elements(8);
    -- CP-element group 125:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1125_entry_sample_req_ps
      -- CP-element group 125: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1125_entry_sample_req
      -- 
    phi_stmt_1125_entry_sample_req_1800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1125_entry_sample_req_1800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(125), ack => phi_stmt_1125_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(125) is bound as output of CP function.
    -- CP-element group 126:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1125_phi_mux_ack_ps
      -- CP-element group 126: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1125_phi_mux_ack
      -- 
    phi_stmt_1125_phi_mux_ack_1803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1125_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(126)); -- 
    -- CP-element group 127:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (4) 
      -- CP-element group 127: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_3_1127_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_3_1127_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_3_1127_sample_completed__ps
      -- CP-element group 127: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_3_1127_sample_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(127) is bound as output of CP function.
    -- CP-element group 128:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_3_1127_update_start_
      -- CP-element group 128: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_3_1127_update_start__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(128) is bound as output of CP function.
    -- CP-element group 129:  join  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	130 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_3_1127_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(129) <= outputPort_3_Daemon_CP_1538_elements(130);
    -- CP-element group 130:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	129 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_3_1127_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(130) is a control-delay.
    cp_element_130_delay: control_delay_element  generic map(name => " 130_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_1538_elements(128), ack => outputPort_3_Daemon_CP_1538_elements(130), clk => clk, reset =>reset);
    -- CP-element group 131:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (4) 
      -- CP-element group 131: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_active_packet_1128_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_active_packet_1128_Sample/req
      -- CP-element group 131: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_active_packet_1128_sample_start__ps
      -- CP-element group 131: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_active_packet_1128_sample_start_
      -- 
    req_1824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(131), ack => next_active_packet_1192_1128_buf_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(131) is bound as output of CP function.
    -- CP-element group 132:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (4) 
      -- CP-element group 132: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_active_packet_1128_update_start_
      -- CP-element group 132: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_active_packet_1128_update_start__ps
      -- CP-element group 132: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_active_packet_1128_Update/req
      -- CP-element group 132: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_active_packet_1128_Update/$entry
      -- 
    req_1829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(132), ack => next_active_packet_1192_1128_buf_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(132) is bound as output of CP function.
    -- CP-element group 133:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_active_packet_1128_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_active_packet_1128_Sample/ack
      -- CP-element group 133: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_active_packet_1128_sample_completed__ps
      -- CP-element group 133: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_active_packet_1128_sample_completed_
      -- 
    ack_1825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_1192_1128_buf_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(133)); -- 
    -- CP-element group 134:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_active_packet_1128_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_active_packet_1128_update_completed__ps
      -- CP-element group 134: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_active_packet_1128_Update/ack
      -- CP-element group 134: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_active_packet_1128_Update/$exit
      -- 
    ack_1830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_1192_1128_buf_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(134)); -- 
    -- CP-element group 135:  join  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	9 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	12 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	11 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1129_sample_start_
      -- 
    outputPort_3_Daemon_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	9 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	155 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	13 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1129_update_start_
      -- 
    outputPort_3_Daemon_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(9) & outputPort_3_Daemon_CP_1538_elements(155);
      gj_outputPort_3_Daemon_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	11 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1129_sample_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(137) <= outputPort_3_Daemon_CP_1538_elements(11);
    -- CP-element group 138:  join  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	12 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1129_sample_completed__ps
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(138) is bound as output of CP function.
    -- CP-element group 139:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	13 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1129_update_start__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(139) <= outputPort_3_Daemon_CP_1538_elements(13);
    -- CP-element group 140:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	154 
    -- CP-element group 140: 	14 
    -- CP-element group 140:  members (2) 
      -- CP-element group 140: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1129_update_completed__ps
      -- CP-element group 140: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1129_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(140) is bound as output of CP function.
    -- CP-element group 141:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	7 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1129_loopback_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(141) <= outputPort_3_Daemon_CP_1538_elements(7);
    -- CP-element group 142:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1129_loopback_sample_req_ps
      -- CP-element group 142: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1129_loopback_sample_req
      -- 
    phi_stmt_1129_loopback_sample_req_1841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1129_loopback_sample_req_1841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(142), ack => phi_stmt_1129_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(142) is bound as output of CP function.
    -- CP-element group 143:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	8 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1129_entry_trigger
      -- 
    outputPort_3_Daemon_CP_1538_elements(143) <= outputPort_3_Daemon_CP_1538_elements(8);
    -- CP-element group 144:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1129_entry_sample_req
      -- CP-element group 144: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1129_entry_sample_req_ps
      -- 
    phi_stmt_1129_entry_sample_req_1844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1129_entry_sample_req_1844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(144), ack => phi_stmt_1129_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1129_phi_mux_ack_ps
      -- CP-element group 145: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/phi_stmt_1129_phi_mux_ack
      -- 
    phi_stmt_1129_phi_mux_ack_1847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1129_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(145)); -- 
    -- CP-element group 146:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (4) 
      -- CP-element group 146: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_3_1131_sample_completed_
      -- CP-element group 146: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_3_1131_sample_start__ps
      -- CP-element group 146: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_3_1131_sample_completed__ps
      -- CP-element group 146: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_3_1131_sample_start_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(146) is bound as output of CP function.
    -- CP-element group 147:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (2) 
      -- CP-element group 147: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_3_1131_update_start__ps
      -- CP-element group 147: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_3_1131_update_start_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(147) is bound as output of CP function.
    -- CP-element group 148:  join  transition  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	149 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (1) 
      -- CP-element group 148: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_3_1131_update_completed__ps
      -- 
    outputPort_3_Daemon_CP_1538_elements(148) <= outputPort_3_Daemon_CP_1538_elements(149);
    -- CP-element group 149:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	148 
    -- CP-element group 149:  members (1) 
      -- CP-element group 149: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_ZERO_3_1131_update_completed_
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(149) is a control-delay.
    cp_element_149_delay: control_delay_element  generic map(name => " 149_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_1538_elements(147), ack => outputPort_3_Daemon_CP_1538_elements(149), clk => clk, reset =>reset);
    -- CP-element group 150:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (4) 
      -- CP-element group 150: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_pkt_priority_1132_sample_start__ps
      -- CP-element group 150: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_pkt_priority_1132_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_pkt_priority_1132_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_pkt_priority_1132_Sample/req
      -- 
    req_1868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(150), ack => next_pkt_priority_1192_1132_buf_req_0); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(150) is bound as output of CP function.
    -- CP-element group 151:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (4) 
      -- CP-element group 151: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_pkt_priority_1132_update_start__ps
      -- CP-element group 151: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_pkt_priority_1132_update_start_
      -- CP-element group 151: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_pkt_priority_1132_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_pkt_priority_1132_Update/req
      -- 
    req_1873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(151), ack => next_pkt_priority_1192_1132_buf_req_1); -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(151) is bound as output of CP function.
    -- CP-element group 152:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (4) 
      -- CP-element group 152: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_pkt_priority_1132_sample_completed__ps
      -- CP-element group 152: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_pkt_priority_1132_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_pkt_priority_1132_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_pkt_priority_1132_Sample/ack
      -- 
    ack_1869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pkt_priority_1192_1132_buf_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(152)); -- 
    -- CP-element group 153:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (4) 
      -- CP-element group 153: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_pkt_priority_1132_update_completed__ps
      -- CP-element group 153: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_pkt_priority_1132_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_pkt_priority_1132_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/R_next_pkt_priority_1132_Update/ack
      -- 
    ack_1874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pkt_priority_1192_1132_buf_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	121 
    -- CP-element group 154: 	102 
    -- CP-element group 154: 	60 
    -- CP-element group 154: 	81 
    -- CP-element group 154: 	140 
    -- CP-element group 154: 	20 
    -- CP-element group 154: 	39 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/WPIPE_out_data_3_1312_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/WPIPE_out_data_3_1312_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/WPIPE_out_data_3_1312_Sample/req
      -- 
    req_1883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(154), ack => WPIPE_out_data_3_1312_inst_req_0); -- 
    outputPort_3_Daemon_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(121) & outputPort_3_Daemon_CP_1538_elements(102) & outputPort_3_Daemon_CP_1538_elements(60) & outputPort_3_Daemon_CP_1538_elements(81) & outputPort_3_Daemon_CP_1538_elements(140) & outputPort_3_Daemon_CP_1538_elements(20) & outputPort_3_Daemon_CP_1538_elements(39) & outputPort_3_Daemon_CP_1538_elements(156);
      gj_outputPort_3_Daemon_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	119 
    -- CP-element group 155: 	136 
    -- CP-element group 155: 	56 
    -- CP-element group 155: 	98 
    -- CP-element group 155: 	77 
    -- CP-element group 155: 	16 
    -- CP-element group 155: 	35 
    -- CP-element group 155:  members (6) 
      -- CP-element group 155: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/WPIPE_out_data_3_1312_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/WPIPE_out_data_3_1312_update_start_
      -- CP-element group 155: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/WPIPE_out_data_3_1312_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/WPIPE_out_data_3_1312_Sample/ack
      -- CP-element group 155: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/WPIPE_out_data_3_1312_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/WPIPE_out_data_3_1312_Update/req
      -- 
    ack_1884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_3_1312_inst_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(155)); -- 
    req_1888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_3_Daemon_CP_1538_elements(155), ack => WPIPE_out_data_3_1312_inst_req_1); -- 
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	154 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/WPIPE_out_data_3_1312_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/WPIPE_out_data_3_1312_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/WPIPE_out_data_3_1312_Update/ack
      -- 
    ack_1889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_3_1312_inst_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(156)); -- 
    -- CP-element group 157:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	9 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	10 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group outputPort_3_Daemon_CP_1538_elements(157) is a control-delay.
    cp_element_157_delay: control_delay_element  generic map(name => " 157_delay", delay_value => 1)  port map(req => outputPort_3_Daemon_CP_1538_elements(9), ack => outputPort_3_Daemon_CP_1538_elements(157), clk => clk, reset =>reset);
    -- CP-element group 158:  join  transition  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: 	12 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	6 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_1098/do_while_stmt_1099/do_while_stmt_1099_loop_body/$exit
      -- 
    outputPort_3_Daemon_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_3_Daemon_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_3_Daemon_CP_1538_elements(156) & outputPort_3_Daemon_CP_1538_elements(12);
      gj_outputPort_3_Daemon_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	5 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (2) 
      -- CP-element group 159: 	 branch_block_stmt_1098/do_while_stmt_1099/loop_exit/$exit
      -- CP-element group 159: 	 branch_block_stmt_1098/do_while_stmt_1099/loop_exit/ack
      -- 
    ack_1894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1099_branch_ack_0, ack => outputPort_3_Daemon_CP_1538_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	5 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (2) 
      -- CP-element group 160: 	 branch_block_stmt_1098/do_while_stmt_1099/loop_taken/$exit
      -- CP-element group 160: 	 branch_block_stmt_1098/do_while_stmt_1099/loop_taken/ack
      -- 
    ack_1898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1099_branch_ack_1, ack => outputPort_3_Daemon_CP_1538_elements(160)); -- 
    -- CP-element group 161:  transition  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	3 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	1 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_1098/do_while_stmt_1099/$exit
      -- 
    outputPort_3_Daemon_CP_1538_elements(161) <= outputPort_3_Daemon_CP_1538_elements(3);
    outputPort_3_Daemon_do_while_stmt_1099_terminator_1899: loop_terminator -- 
      generic map (name => " outputPort_3_Daemon_do_while_stmt_1099_terminator_1899", max_iterations_in_flight =>7) 
      port map(loop_body_exit => outputPort_3_Daemon_CP_1538_elements(6),loop_continue => outputPort_3_Daemon_CP_1538_elements(160),loop_terminate => outputPort_3_Daemon_CP_1538_elements(159),loop_back => outputPort_3_Daemon_CP_1538_elements(4),loop_exit => outputPort_3_Daemon_CP_1538_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1101_phi_seq_1611_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_1538_elements(23);
      outputPort_3_Daemon_CP_1538_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(26);
      outputPort_3_Daemon_CP_1538_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(28);
      outputPort_3_Daemon_CP_1538_elements(24) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_1538_elements(21);
      outputPort_3_Daemon_CP_1538_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(32);
      outputPort_3_Daemon_CP_1538_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(33);
      outputPort_3_Daemon_CP_1538_elements(22) <= phi_mux_reqs(1);
      phi_stmt_1101_phi_seq_1611 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1101_phi_seq_1611") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_1538_elements(17), 
          phi_sample_ack => outputPort_3_Daemon_CP_1538_elements(18), 
          phi_update_req => outputPort_3_Daemon_CP_1538_elements(19), 
          phi_update_ack => outputPort_3_Daemon_CP_1538_elements(20), 
          phi_mux_ack => outputPort_3_Daemon_CP_1538_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1105_phi_seq_1655_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_1538_elements(42);
      outputPort_3_Daemon_CP_1538_elements(45)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(45);
      outputPort_3_Daemon_CP_1538_elements(46)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(47);
      outputPort_3_Daemon_CP_1538_elements(43) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_1538_elements(40);
      outputPort_3_Daemon_CP_1538_elements(49)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(53);
      outputPort_3_Daemon_CP_1538_elements(50)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(54);
      outputPort_3_Daemon_CP_1538_elements(41) <= phi_mux_reqs(1);
      phi_stmt_1105_phi_seq_1655 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1105_phi_seq_1655") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_1538_elements(36), 
          phi_sample_ack => outputPort_3_Daemon_CP_1538_elements(37), 
          phi_update_req => outputPort_3_Daemon_CP_1538_elements(38), 
          phi_update_ack => outputPort_3_Daemon_CP_1538_elements(39), 
          phi_mux_ack => outputPort_3_Daemon_CP_1538_elements(44), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1110_phi_seq_1699_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_1538_elements(63);
      outputPort_3_Daemon_CP_1538_elements(66)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(66);
      outputPort_3_Daemon_CP_1538_elements(67)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(68);
      outputPort_3_Daemon_CP_1538_elements(64) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_1538_elements(61);
      outputPort_3_Daemon_CP_1538_elements(70)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(74);
      outputPort_3_Daemon_CP_1538_elements(71)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(75);
      outputPort_3_Daemon_CP_1538_elements(62) <= phi_mux_reqs(1);
      phi_stmt_1110_phi_seq_1699 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1110_phi_seq_1699") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_1538_elements(57), 
          phi_sample_ack => outputPort_3_Daemon_CP_1538_elements(58), 
          phi_update_req => outputPort_3_Daemon_CP_1538_elements(59), 
          phi_update_ack => outputPort_3_Daemon_CP_1538_elements(60), 
          phi_mux_ack => outputPort_3_Daemon_CP_1538_elements(65), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1115_phi_seq_1743_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_1538_elements(84);
      outputPort_3_Daemon_CP_1538_elements(87)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(87);
      outputPort_3_Daemon_CP_1538_elements(88)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(89);
      outputPort_3_Daemon_CP_1538_elements(85) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_1538_elements(82);
      outputPort_3_Daemon_CP_1538_elements(91)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(95);
      outputPort_3_Daemon_CP_1538_elements(92)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(96);
      outputPort_3_Daemon_CP_1538_elements(83) <= phi_mux_reqs(1);
      phi_stmt_1115_phi_seq_1743 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1115_phi_seq_1743") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_1538_elements(78), 
          phi_sample_ack => outputPort_3_Daemon_CP_1538_elements(79), 
          phi_update_req => outputPort_3_Daemon_CP_1538_elements(80), 
          phi_update_ack => outputPort_3_Daemon_CP_1538_elements(81), 
          phi_mux_ack => outputPort_3_Daemon_CP_1538_elements(86), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1120_phi_seq_1787_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_1538_elements(105);
      outputPort_3_Daemon_CP_1538_elements(108)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(108);
      outputPort_3_Daemon_CP_1538_elements(109)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(110);
      outputPort_3_Daemon_CP_1538_elements(106) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_1538_elements(103);
      outputPort_3_Daemon_CP_1538_elements(112)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(116);
      outputPort_3_Daemon_CP_1538_elements(113)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(117);
      outputPort_3_Daemon_CP_1538_elements(104) <= phi_mux_reqs(1);
      phi_stmt_1120_phi_seq_1787 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1120_phi_seq_1787") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_1538_elements(99), 
          phi_sample_ack => outputPort_3_Daemon_CP_1538_elements(100), 
          phi_update_req => outputPort_3_Daemon_CP_1538_elements(101), 
          phi_update_ack => outputPort_3_Daemon_CP_1538_elements(102), 
          phi_mux_ack => outputPort_3_Daemon_CP_1538_elements(107), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1125_phi_seq_1831_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_1538_elements(124);
      outputPort_3_Daemon_CP_1538_elements(127)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(127);
      outputPort_3_Daemon_CP_1538_elements(128)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(129);
      outputPort_3_Daemon_CP_1538_elements(125) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_1538_elements(122);
      outputPort_3_Daemon_CP_1538_elements(131)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(133);
      outputPort_3_Daemon_CP_1538_elements(132)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(134);
      outputPort_3_Daemon_CP_1538_elements(123) <= phi_mux_reqs(1);
      phi_stmt_1125_phi_seq_1831 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1125_phi_seq_1831") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_1538_elements(11), 
          phi_sample_ack => outputPort_3_Daemon_CP_1538_elements(120), 
          phi_update_req => outputPort_3_Daemon_CP_1538_elements(13), 
          phi_update_ack => outputPort_3_Daemon_CP_1538_elements(121), 
          phi_mux_ack => outputPort_3_Daemon_CP_1538_elements(126), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1129_phi_seq_1875_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_3_Daemon_CP_1538_elements(143);
      outputPort_3_Daemon_CP_1538_elements(146)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(146);
      outputPort_3_Daemon_CP_1538_elements(147)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_3_Daemon_CP_1538_elements(148);
      outputPort_3_Daemon_CP_1538_elements(144) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_3_Daemon_CP_1538_elements(141);
      outputPort_3_Daemon_CP_1538_elements(150)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(152);
      outputPort_3_Daemon_CP_1538_elements(151)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_3_Daemon_CP_1538_elements(153);
      outputPort_3_Daemon_CP_1538_elements(142) <= phi_mux_reqs(1);
      phi_stmt_1129_phi_seq_1875 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1129_phi_seq_1875") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_3_Daemon_CP_1538_elements(137), 
          phi_sample_ack => outputPort_3_Daemon_CP_1538_elements(138), 
          phi_update_req => outputPort_3_Daemon_CP_1538_elements(139), 
          phi_update_ack => outputPort_3_Daemon_CP_1538_elements(140), 
          phi_mux_ack => outputPort_3_Daemon_CP_1538_elements(145), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1563_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= outputPort_3_Daemon_CP_1538_elements(7);
        preds(1)  <= outputPort_3_Daemon_CP_1538_elements(8);
        entry_tmerge_1563 : transition_merge -- 
          generic map(name => " entry_tmerge_1563")
          port map (preds => preds, symbol_out => outputPort_3_Daemon_CP_1538_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u3_u1_1157_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1163_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1170_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1176_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1222_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1230_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1238_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1246_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1252_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1259_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1267_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1274_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1285_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1291_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1298_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1304_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_1203_wire : std_logic_vector(0 downto 0);
    signal MUX_1160_wire : std_logic_vector(0 downto 0);
    signal MUX_1166_wire : std_logic_vector(0 downto 0);
    signal MUX_1173_wire : std_logic_vector(0 downto 0);
    signal MUX_1179_wire : std_logic_vector(0 downto 0);
    signal MUX_1214_wire : std_logic_vector(7 downto 0);
    signal MUX_1256_wire : std_logic_vector(31 downto 0);
    signal MUX_1263_wire : std_logic_vector(31 downto 0);
    signal MUX_1271_wire : std_logic_vector(31 downto 0);
    signal MUX_1278_wire : std_logic_vector(31 downto 0);
    signal MUX_1288_wire : std_logic_vector(0 downto 0);
    signal MUX_1294_wire : std_logic_vector(0 downto 0);
    signal MUX_1301_wire : std_logic_vector(0 downto 0);
    signal MUX_1307_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1219_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1227_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1235_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1243_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1167_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1180_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1196_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1199_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1200_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1295_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1308_wire : std_logic_vector(0 downto 0);
    signal OR_u32_u32_1264_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_1279_wire : std_logic_vector(31 downto 0);
    signal RPIPE_noblock_obuf_1_3_1109_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_2_3_1114_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_3_3_1119_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_4_3_1124_wire : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1107_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1112_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1117_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1122_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_3_1127_wire_constant : std_logic_vector(2 downto 0);
    signal R_ZERO_3_1131_wire_constant : std_logic_vector(2 downto 0);
    signal R_ZERO_8_1103_wire_constant : std_logic_vector(7 downto 0);
    signal SUB_u8_u8_1212_wire : std_logic_vector(7 downto 0);
    signal active_packet_1125 : std_logic_vector(2 downto 0);
    signal data_to_out_1281 : std_logic_vector(31 downto 0);
    signal down_counter_1101 : std_logic_vector(7 downto 0);
    signal konst_1136_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1141_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1146_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1151_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1156_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1159_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1162_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1165_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1169_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1172_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1175_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1178_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1202_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1208_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1211_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1221_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1229_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1237_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1245_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1251_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1255_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1258_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1262_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1266_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1270_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1273_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1277_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1284_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1287_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1290_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1293_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1297_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1300_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1303_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1306_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1316_wire_constant : std_logic_vector(0 downto 0);
    signal next_active_packet_1192 : std_logic_vector(2 downto 0);
    signal next_active_packet_1192_1128_buffered : std_logic_vector(2 downto 0);
    signal next_down_counter_1216 : std_logic_vector(7 downto 0);
    signal next_down_counter_1216_1104_buffered : std_logic_vector(7 downto 0);
    signal next_pkt_priority_1192 : std_logic_vector(2 downto 0);
    signal next_pkt_priority_1192_1132_buffered : std_logic_vector(2 downto 0);
    signal p1_valid_1138 : std_logic_vector(0 downto 0);
    signal p2_valid_1143 : std_logic_vector(0 downto 0);
    signal p3_valid_1148 : std_logic_vector(0 downto 0);
    signal p4_valid_1153 : std_logic_vector(0 downto 0);
    signal pkt_1_e_word_1105 : std_logic_vector(32 downto 0);
    signal pkt_2_e_word_1110 : std_logic_vector(32 downto 0);
    signal pkt_3_e_word_1115 : std_logic_vector(32 downto 0);
    signal pkt_4_e_word_1120 : std_logic_vector(32 downto 0);
    signal pkt_priority_1129 : std_logic_vector(2 downto 0);
    signal read_from_1_1224 : std_logic_vector(0 downto 0);
    signal read_from_2_1232 : std_logic_vector(0 downto 0);
    signal read_from_3_1240 : std_logic_vector(0 downto 0);
    signal read_from_4_1248 : std_logic_vector(0 downto 0);
    signal send_flag_1310 : std_logic_vector(0 downto 0);
    signal slice_1254_wire : std_logic_vector(31 downto 0);
    signal slice_1261_wire : std_logic_vector(31 downto 0);
    signal slice_1269_wire : std_logic_vector(31 downto 0);
    signal slice_1276_wire : std_logic_vector(31 downto 0);
    signal started_new_packet_1205 : std_logic_vector(0 downto 0);
    signal valid_active_pkt_word_read_1182 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_ZERO_33_1107_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1112_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1117_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1122_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_3_1127_wire_constant <= "000";
    R_ZERO_3_1131_wire_constant <= "000";
    R_ZERO_8_1103_wire_constant <= "00000000";
    konst_1136_wire_constant <= "000000000000000000000000000100000";
    konst_1141_wire_constant <= "000000000000000000000000000100000";
    konst_1146_wire_constant <= "000000000000000000000000000100000";
    konst_1151_wire_constant <= "000000000000000000000000000100000";
    konst_1156_wire_constant <= "001";
    konst_1159_wire_constant <= "0";
    konst_1162_wire_constant <= "010";
    konst_1165_wire_constant <= "0";
    konst_1169_wire_constant <= "011";
    konst_1172_wire_constant <= "0";
    konst_1175_wire_constant <= "100";
    konst_1178_wire_constant <= "0";
    konst_1202_wire_constant <= "00000000";
    konst_1208_wire_constant <= "00111111";
    konst_1211_wire_constant <= "00000001";
    konst_1221_wire_constant <= "001";
    konst_1229_wire_constant <= "010";
    konst_1237_wire_constant <= "011";
    konst_1245_wire_constant <= "100";
    konst_1251_wire_constant <= "001";
    konst_1255_wire_constant <= "00000000000000000000000000000000";
    konst_1258_wire_constant <= "010";
    konst_1262_wire_constant <= "00000000000000000000000000000000";
    konst_1266_wire_constant <= "011";
    konst_1270_wire_constant <= "00000000000000000000000000000000";
    konst_1273_wire_constant <= "100";
    konst_1277_wire_constant <= "00000000000000000000000000000000";
    konst_1284_wire_constant <= "001";
    konst_1287_wire_constant <= "0";
    konst_1290_wire_constant <= "010";
    konst_1293_wire_constant <= "0";
    konst_1297_wire_constant <= "011";
    konst_1300_wire_constant <= "0";
    konst_1303_wire_constant <= "100";
    konst_1306_wire_constant <= "0";
    konst_1316_wire_constant <= "1";
    phi_stmt_1101: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_8_1103_wire_constant & next_down_counter_1216_1104_buffered;
      req <= phi_stmt_1101_req_0 & phi_stmt_1101_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1101",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1101_ack_0,
          idata => idata,
          odata => down_counter_1101,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1101
    phi_stmt_1105: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1107_wire_constant & RPIPE_noblock_obuf_1_3_1109_wire;
      req <= phi_stmt_1105_req_0 & phi_stmt_1105_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1105",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1105_ack_0,
          idata => idata,
          odata => pkt_1_e_word_1105,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1105
    phi_stmt_1110: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1112_wire_constant & RPIPE_noblock_obuf_2_3_1114_wire;
      req <= phi_stmt_1110_req_0 & phi_stmt_1110_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1110",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1110_ack_0,
          idata => idata,
          odata => pkt_2_e_word_1110,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1110
    phi_stmt_1115: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1117_wire_constant & RPIPE_noblock_obuf_3_3_1119_wire;
      req <= phi_stmt_1115_req_0 & phi_stmt_1115_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1115",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1115_ack_0,
          idata => idata,
          odata => pkt_3_e_word_1115,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1115
    phi_stmt_1120: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1122_wire_constant & RPIPE_noblock_obuf_4_3_1124_wire;
      req <= phi_stmt_1120_req_0 & phi_stmt_1120_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1120",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1120_ack_0,
          idata => idata,
          odata => pkt_4_e_word_1120,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1120
    phi_stmt_1125: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_3_1127_wire_constant & next_active_packet_1192_1128_buffered;
      req <= phi_stmt_1125_req_0 & phi_stmt_1125_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1125",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1125_ack_0,
          idata => idata,
          odata => active_packet_1125,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1125
    phi_stmt_1129: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_3_1131_wire_constant & next_pkt_priority_1192_1132_buffered;
      req <= phi_stmt_1129_req_0 & phi_stmt_1129_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1129",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1129_ack_0,
          idata => idata,
          odata => pkt_priority_1129,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1129
    -- flow-through select operator MUX_1160_inst
    MUX_1160_wire <= p1_valid_1138 when (EQ_u3_u1_1157_wire(0) /=  '0') else konst_1159_wire_constant;
    -- flow-through select operator MUX_1166_inst
    MUX_1166_wire <= p2_valid_1143 when (EQ_u3_u1_1163_wire(0) /=  '0') else konst_1165_wire_constant;
    -- flow-through select operator MUX_1173_inst
    MUX_1173_wire <= p3_valid_1148 when (EQ_u3_u1_1170_wire(0) /=  '0') else konst_1172_wire_constant;
    -- flow-through select operator MUX_1179_inst
    MUX_1179_wire <= p4_valid_1153 when (EQ_u3_u1_1176_wire(0) /=  '0') else konst_1178_wire_constant;
    -- flow-through select operator MUX_1214_inst
    MUX_1214_wire <= SUB_u8_u8_1212_wire when (valid_active_pkt_word_read_1182(0) /=  '0') else down_counter_1101;
    -- flow-through select operator MUX_1215_inst
    next_down_counter_1216 <= konst_1208_wire_constant when (started_new_packet_1205(0) /=  '0') else MUX_1214_wire;
    -- flow-through select operator MUX_1256_inst
    MUX_1256_wire <= slice_1254_wire when (EQ_u3_u1_1252_wire(0) /=  '0') else konst_1255_wire_constant;
    -- flow-through select operator MUX_1263_inst
    MUX_1263_wire <= slice_1261_wire when (EQ_u3_u1_1259_wire(0) /=  '0') else konst_1262_wire_constant;
    -- flow-through select operator MUX_1271_inst
    MUX_1271_wire <= slice_1269_wire when (EQ_u3_u1_1267_wire(0) /=  '0') else konst_1270_wire_constant;
    -- flow-through select operator MUX_1278_inst
    MUX_1278_wire <= slice_1276_wire when (EQ_u3_u1_1274_wire(0) /=  '0') else konst_1277_wire_constant;
    -- flow-through select operator MUX_1288_inst
    MUX_1288_wire <= p1_valid_1138 when (EQ_u3_u1_1285_wire(0) /=  '0') else konst_1287_wire_constant;
    -- flow-through select operator MUX_1294_inst
    MUX_1294_wire <= p2_valid_1143 when (EQ_u3_u1_1291_wire(0) /=  '0') else konst_1293_wire_constant;
    -- flow-through select operator MUX_1301_inst
    MUX_1301_wire <= p3_valid_1148 when (EQ_u3_u1_1298_wire(0) /=  '0') else konst_1300_wire_constant;
    -- flow-through select operator MUX_1307_inst
    MUX_1307_wire <= p4_valid_1153 when (EQ_u3_u1_1304_wire(0) /=  '0') else konst_1306_wire_constant;
    -- flow-through slice operator slice_1254_inst
    slice_1254_wire <= pkt_1_e_word_1105(31 downto 0);
    -- flow-through slice operator slice_1261_inst
    slice_1261_wire <= pkt_2_e_word_1110(31 downto 0);
    -- flow-through slice operator slice_1269_inst
    slice_1269_wire <= pkt_3_e_word_1115(31 downto 0);
    -- flow-through slice operator slice_1276_inst
    slice_1276_wire <= pkt_4_e_word_1120(31 downto 0);
    next_active_packet_1192_1128_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_active_packet_1192_1128_buf_req_0;
      next_active_packet_1192_1128_buf_ack_0<= wack(0);
      rreq(0) <= next_active_packet_1192_1128_buf_req_1;
      next_active_packet_1192_1128_buf_ack_1<= rack(0);
      next_active_packet_1192_1128_buf : InterlockBuffer generic map ( -- 
        name => "next_active_packet_1192_1128_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_active_packet_1192,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_active_packet_1192_1128_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_down_counter_1216_1104_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_down_counter_1216_1104_buf_req_0;
      next_down_counter_1216_1104_buf_ack_0<= wack(0);
      rreq(0) <= next_down_counter_1216_1104_buf_req_1;
      next_down_counter_1216_1104_buf_ack_1<= rack(0);
      next_down_counter_1216_1104_buf : InterlockBuffer generic map ( -- 
        name => "next_down_counter_1216_1104_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_down_counter_1216,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_down_counter_1216_1104_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_pkt_priority_1192_1132_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_pkt_priority_1192_1132_buf_req_0;
      next_pkt_priority_1192_1132_buf_ack_0<= wack(0);
      rreq(0) <= next_pkt_priority_1192_1132_buf_req_1;
      next_pkt_priority_1192_1132_buf_ack_1<= rack(0);
      next_pkt_priority_1192_1132_buf : InterlockBuffer generic map ( -- 
        name => "next_pkt_priority_1192_1132_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_pkt_priority_1192,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_pkt_priority_1192_1132_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1099_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1316_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1099_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1099_branch_req_0,
          ack0 => do_while_stmt_1099_branch_ack_0,
          ack1 => do_while_stmt_1099_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator AND_u1_u1_1204_inst
    process(OR_u1_u1_1200_wire, EQ_u8_u1_1203_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(OR_u1_u1_1200_wire, EQ_u8_u1_1203_wire, tmp_var);
      started_new_packet_1205 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_1137_inst
    process(pkt_1_e_word_1105) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_1_e_word_1105, konst_1136_wire_constant, tmp_var);
      p1_valid_1138 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_1142_inst
    process(pkt_2_e_word_1110) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_2_e_word_1110, konst_1141_wire_constant, tmp_var);
      p2_valid_1143 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_1147_inst
    process(pkt_3_e_word_1115) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_3_e_word_1115, konst_1146_wire_constant, tmp_var);
      p3_valid_1148 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_1152_inst
    process(pkt_4_e_word_1120) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_4_e_word_1120, konst_1151_wire_constant, tmp_var);
      p4_valid_1153 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1157_inst
    process(active_packet_1125) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1125, konst_1156_wire_constant, tmp_var);
      EQ_u3_u1_1157_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1163_inst
    process(active_packet_1125) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1125, konst_1162_wire_constant, tmp_var);
      EQ_u3_u1_1163_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1170_inst
    process(active_packet_1125) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1125, konst_1169_wire_constant, tmp_var);
      EQ_u3_u1_1170_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1176_inst
    process(active_packet_1125) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1125, konst_1175_wire_constant, tmp_var);
      EQ_u3_u1_1176_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1222_inst
    process(next_active_packet_1192) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1192, konst_1221_wire_constant, tmp_var);
      EQ_u3_u1_1222_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1230_inst
    process(next_active_packet_1192) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1192, konst_1229_wire_constant, tmp_var);
      EQ_u3_u1_1230_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1238_inst
    process(next_active_packet_1192) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1192, konst_1237_wire_constant, tmp_var);
      EQ_u3_u1_1238_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1246_inst
    process(next_active_packet_1192) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1192, konst_1245_wire_constant, tmp_var);
      EQ_u3_u1_1246_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1252_inst
    process(next_active_packet_1192) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1192, konst_1251_wire_constant, tmp_var);
      EQ_u3_u1_1252_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1259_inst
    process(next_active_packet_1192) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1192, konst_1258_wire_constant, tmp_var);
      EQ_u3_u1_1259_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1267_inst
    process(next_active_packet_1192) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1192, konst_1266_wire_constant, tmp_var);
      EQ_u3_u1_1267_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1274_inst
    process(next_active_packet_1192) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1192, konst_1273_wire_constant, tmp_var);
      EQ_u3_u1_1274_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1285_inst
    process(next_active_packet_1192) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1192, konst_1284_wire_constant, tmp_var);
      EQ_u3_u1_1285_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1291_inst
    process(next_active_packet_1192) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1192, konst_1290_wire_constant, tmp_var);
      EQ_u3_u1_1291_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1298_inst
    process(next_active_packet_1192) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1192, konst_1297_wire_constant, tmp_var);
      EQ_u3_u1_1298_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1304_inst
    process(next_active_packet_1192) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1192, konst_1303_wire_constant, tmp_var);
      EQ_u3_u1_1304_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_1203_inst
    process(down_counter_1101) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(down_counter_1101, konst_1202_wire_constant, tmp_var);
      EQ_u8_u1_1203_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1219_inst
    process(p1_valid_1138) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_1138, tmp_var);
      NOT_u1_u1_1219_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1227_inst
    process(p2_valid_1143) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_1143, tmp_var);
      NOT_u1_u1_1227_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1235_inst
    process(p3_valid_1148) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_1148, tmp_var);
      NOT_u1_u1_1235_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1243_inst
    process(p4_valid_1153) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_1153, tmp_var);
      NOT_u1_u1_1243_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1167_inst
    process(MUX_1160_wire, MUX_1166_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1160_wire, MUX_1166_wire, tmp_var);
      OR_u1_u1_1167_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1180_inst
    process(MUX_1173_wire, MUX_1179_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1173_wire, MUX_1179_wire, tmp_var);
      OR_u1_u1_1180_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1181_inst
    process(OR_u1_u1_1167_wire, OR_u1_u1_1180_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1167_wire, OR_u1_u1_1180_wire, tmp_var);
      valid_active_pkt_word_read_1182 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1196_inst
    process(p1_valid_1138, p2_valid_1143) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(p1_valid_1138, p2_valid_1143, tmp_var);
      OR_u1_u1_1196_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1199_inst
    process(p3_valid_1148, p4_valid_1153) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(p3_valid_1148, p4_valid_1153, tmp_var);
      OR_u1_u1_1199_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1200_inst
    process(OR_u1_u1_1196_wire, OR_u1_u1_1199_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1196_wire, OR_u1_u1_1199_wire, tmp_var);
      OR_u1_u1_1200_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1223_inst
    process(NOT_u1_u1_1219_wire, EQ_u3_u1_1222_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1219_wire, EQ_u3_u1_1222_wire, tmp_var);
      read_from_1_1224 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1231_inst
    process(NOT_u1_u1_1227_wire, EQ_u3_u1_1230_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1227_wire, EQ_u3_u1_1230_wire, tmp_var);
      read_from_2_1232 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1239_inst
    process(NOT_u1_u1_1235_wire, EQ_u3_u1_1238_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1235_wire, EQ_u3_u1_1238_wire, tmp_var);
      read_from_3_1240 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1247_inst
    process(NOT_u1_u1_1243_wire, EQ_u3_u1_1246_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1243_wire, EQ_u3_u1_1246_wire, tmp_var);
      read_from_4_1248 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1295_inst
    process(MUX_1288_wire, MUX_1294_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1288_wire, MUX_1294_wire, tmp_var);
      OR_u1_u1_1295_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1308_inst
    process(MUX_1301_wire, MUX_1307_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1301_wire, MUX_1307_wire, tmp_var);
      OR_u1_u1_1308_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1309_inst
    process(OR_u1_u1_1295_wire, OR_u1_u1_1308_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1295_wire, OR_u1_u1_1308_wire, tmp_var);
      send_flag_1310 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1264_inst
    process(MUX_1256_wire, MUX_1263_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1256_wire, MUX_1263_wire, tmp_var);
      OR_u32_u32_1264_wire <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1279_inst
    process(MUX_1271_wire, MUX_1278_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1271_wire, MUX_1278_wire, tmp_var);
      OR_u32_u32_1279_wire <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1280_inst
    process(OR_u32_u32_1264_wire, OR_u32_u32_1279_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u32_u32_1264_wire, OR_u32_u32_1279_wire, tmp_var);
      data_to_out_1281 <= tmp_var; --
    end process;
    -- binary operator SUB_u8_u8_1212_inst
    process(down_counter_1101) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSub_proc(down_counter_1101, konst_1211_wire_constant, tmp_var);
      SUB_u8_u8_1212_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_noblock_obuf_1_3_1109_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_1_3_1109_inst_req_0;
      RPIPE_noblock_obuf_1_3_1109_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_1_3_1109_inst_req_1;
      RPIPE_noblock_obuf_1_3_1109_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_1_1224(0);
      RPIPE_noblock_obuf_1_3_1109_wire <= data_out(32 downto 0);
      noblock_obuf_1_3_read_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_3_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_3_read_0: InputPortRevised -- 
        generic map ( name => "noblock_obuf_1_3_read_0", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_1_3_pipe_read_req(0),
          oack => noblock_obuf_1_3_pipe_read_ack(0),
          odata => noblock_obuf_1_3_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_noblock_obuf_2_3_1114_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_2_3_1114_inst_req_0;
      RPIPE_noblock_obuf_2_3_1114_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_2_3_1114_inst_req_1;
      RPIPE_noblock_obuf_2_3_1114_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_2_1232(0);
      RPIPE_noblock_obuf_2_3_1114_wire <= data_out(32 downto 0);
      noblock_obuf_2_3_read_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_3_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_3_read_1: InputPortRevised -- 
        generic map ( name => "noblock_obuf_2_3_read_1", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_2_3_pipe_read_req(0),
          oack => noblock_obuf_2_3_pipe_read_ack(0),
          odata => noblock_obuf_2_3_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_noblock_obuf_3_3_1119_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_3_3_1119_inst_req_0;
      RPIPE_noblock_obuf_3_3_1119_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_3_3_1119_inst_req_1;
      RPIPE_noblock_obuf_3_3_1119_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_3_1240(0);
      RPIPE_noblock_obuf_3_3_1119_wire <= data_out(32 downto 0);
      noblock_obuf_3_3_read_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_3_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_3_read_2: InputPortRevised -- 
        generic map ( name => "noblock_obuf_3_3_read_2", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_3_3_pipe_read_req(0),
          oack => noblock_obuf_3_3_pipe_read_ack(0),
          odata => noblock_obuf_3_3_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_noblock_obuf_4_3_1124_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_4_3_1124_inst_req_0;
      RPIPE_noblock_obuf_4_3_1124_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_4_3_1124_inst_req_1;
      RPIPE_noblock_obuf_4_3_1124_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_4_1248(0);
      RPIPE_noblock_obuf_4_3_1124_wire <= data_out(32 downto 0);
      noblock_obuf_4_3_read_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_3_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_3_read_3: InputPortRevised -- 
        generic map ( name => "noblock_obuf_4_3_read_3", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_4_3_pipe_read_req(0),
          oack => noblock_obuf_4_3_pipe_read_ack(0),
          odata => noblock_obuf_4_3_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_out_data_3_1312_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_out_data_3_1312_inst_req_0;
      WPIPE_out_data_3_1312_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_out_data_3_1312_inst_req_1;
      WPIPE_out_data_3_1312_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_flag_1310(0);
      data_in <= data_to_out_1281;
      out_data_3_write_0_gI: SplitGuardInterface generic map(name => "out_data_3_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      out_data_3_write_0: OutputPortRevised -- 
        generic map ( name => "out_data_3", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => out_data_3_pipe_write_req(0),
          oack => out_data_3_pipe_write_ack(0),
          odata => out_data_3_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    volatile_operator_prioritySelect_3180: prioritySelect_Volatile port map(down_counter => down_counter_1101, active_packet => active_packet_1125, pkt_priority => pkt_priority_1129, p1_valid => p1_valid_1138, p2_valid => p2_valid_1143, p3_valid => p3_valid_1148, p4_valid => p4_valid_1153, next_active_packet => next_active_packet_1192, next_pkt_priority => next_pkt_priority_1192); 
    -- 
  end Block; -- data_path
  -- 
end outputPort_3_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity outputPort_4_Daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    noblock_obuf_1_4_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_1_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_1_4_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_3_4_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_3_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_3_4_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_2_4_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_2_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_2_4_pipe_read_data : in   std_logic_vector(32 downto 0);
    noblock_obuf_4_4_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_obuf_4_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_obuf_4_4_pipe_read_data : in   std_logic_vector(32 downto 0);
    out_data_4_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_4_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity outputPort_4_Daemon;
architecture outputPort_4_Daemon_arch of outputPort_4_Daemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal outputPort_4_Daemon_CP_1900_start: Boolean;
  signal outputPort_4_Daemon_CP_1900_symbol: Boolean;
  -- volatile/operator module components. 
  component prioritySelect_Volatile is -- 
    port ( -- 
      down_counter : in  std_logic_vector(7 downto 0);
      active_packet : in  std_logic_vector(2 downto 0);
      pkt_priority : in  std_logic_vector(2 downto 0);
      p1_valid : in  std_logic_vector(0 downto 0);
      p2_valid : in  std_logic_vector(0 downto 0);
      p3_valid : in  std_logic_vector(0 downto 0);
      p4_valid : in  std_logic_vector(0 downto 0);
      next_active_packet : out  std_logic_vector(2 downto 0);
      next_pkt_priority : out  std_logic_vector(2 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal RPIPE_noblock_obuf_1_4_1331_inst_ack_1 : boolean;
  signal RPIPE_noblock_obuf_2_4_1336_inst_ack_1 : boolean;
  signal next_down_counter_1438_1326_buf_ack_0 : boolean;
  signal phi_stmt_1337_req_1 : boolean;
  signal RPIPE_noblock_obuf_2_4_1336_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_3_4_1341_inst_ack_1 : boolean;
  signal phi_stmt_1332_req_0 : boolean;
  signal RPIPE_noblock_obuf_3_4_1341_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_2_4_1336_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_1_4_1331_inst_req_1 : boolean;
  signal phi_stmt_1327_ack_0 : boolean;
  signal RPIPE_noblock_obuf_2_4_1336_inst_req_0 : boolean;
  signal phi_stmt_1327_req_1 : boolean;
  signal RPIPE_noblock_obuf_1_4_1331_inst_req_0 : boolean;
  signal phi_stmt_1327_req_0 : boolean;
  signal next_down_counter_1438_1326_buf_req_0 : boolean;
  signal RPIPE_noblock_obuf_1_4_1331_inst_ack_0 : boolean;
  signal phi_stmt_1332_ack_0 : boolean;
  signal phi_stmt_1332_req_1 : boolean;
  signal phi_stmt_1337_req_0 : boolean;
  signal phi_stmt_1337_ack_0 : boolean;
  signal phi_stmt_1323_ack_0 : boolean;
  signal next_down_counter_1438_1326_buf_ack_1 : boolean;
  signal next_down_counter_1438_1326_buf_req_1 : boolean;
  signal do_while_stmt_1321_branch_req_0 : boolean;
  signal phi_stmt_1323_req_0 : boolean;
  signal phi_stmt_1323_req_1 : boolean;
  signal RPIPE_noblock_obuf_4_4_1346_inst_req_1 : boolean;
  signal RPIPE_noblock_obuf_4_4_1346_inst_ack_1 : boolean;
  signal RPIPE_noblock_obuf_4_4_1346_inst_req_0 : boolean;
  signal RPIPE_noblock_obuf_4_4_1346_inst_ack_0 : boolean;
  signal phi_stmt_1342_ack_0 : boolean;
  signal phi_stmt_1342_req_0 : boolean;
  signal phi_stmt_1342_req_1 : boolean;
  signal RPIPE_noblock_obuf_3_4_1341_inst_ack_0 : boolean;
  signal RPIPE_noblock_obuf_3_4_1341_inst_req_0 : boolean;
  signal phi_stmt_1347_req_1 : boolean;
  signal phi_stmt_1347_req_0 : boolean;
  signal phi_stmt_1347_ack_0 : boolean;
  signal next_active_packet_1414_1350_buf_req_0 : boolean;
  signal next_active_packet_1414_1350_buf_ack_0 : boolean;
  signal next_active_packet_1414_1350_buf_req_1 : boolean;
  signal next_active_packet_1414_1350_buf_ack_1 : boolean;
  signal phi_stmt_1351_req_1 : boolean;
  signal phi_stmt_1351_req_0 : boolean;
  signal phi_stmt_1351_ack_0 : boolean;
  signal next_pkt_priority_1414_1354_buf_req_0 : boolean;
  signal next_pkt_priority_1414_1354_buf_ack_0 : boolean;
  signal next_pkt_priority_1414_1354_buf_req_1 : boolean;
  signal next_pkt_priority_1414_1354_buf_ack_1 : boolean;
  signal WPIPE_out_data_4_1534_inst_req_0 : boolean;
  signal WPIPE_out_data_4_1534_inst_ack_0 : boolean;
  signal WPIPE_out_data_4_1534_inst_req_1 : boolean;
  signal WPIPE_out_data_4_1534_inst_ack_1 : boolean;
  signal do_while_stmt_1321_branch_ack_0 : boolean;
  signal do_while_stmt_1321_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "outputPort_4_Daemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  outputPort_4_Daemon_CP_1900_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "outputPort_4_Daemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_4_Daemon_CP_1900_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= outputPort_4_Daemon_CP_1900_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= outputPort_4_Daemon_CP_1900_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  outputPort_4_Daemon_CP_1900: Block -- control-path 
    signal outputPort_4_Daemon_CP_1900_elements: BooleanArray(161 downto 0);
    -- 
  begin -- 
    outputPort_4_Daemon_CP_1900_elements(0) <= outputPort_4_Daemon_CP_1900_start;
    outputPort_4_Daemon_CP_1900_symbol <= outputPort_4_Daemon_CP_1900_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1320/do_while_stmt_1321__entry__
      -- CP-element group 0: 	 branch_block_stmt_1320/$entry
      -- CP-element group 0: 	 branch_block_stmt_1320/branch_block_stmt_1320__entry__
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	161 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1320/do_while_stmt_1321__exit__
      -- CP-element group 1: 	 branch_block_stmt_1320/branch_block_stmt_1320__exit__
      -- CP-element group 1: 	 branch_block_stmt_1320/$exit
      -- CP-element group 1: 	 $exit
      -- 
    outputPort_4_Daemon_CP_1900_elements(1) <= outputPort_4_Daemon_CP_1900_elements(161);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1320/do_while_stmt_1321/$entry
      -- CP-element group 2: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321__entry__
      -- 
    outputPort_4_Daemon_CP_1900_elements(2) <= outputPort_4_Daemon_CP_1900_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	161 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321__exit__
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1320/do_while_stmt_1321/loop_back
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	159 
    -- CP-element group 5: 	160 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1320/do_while_stmt_1321/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1320/do_while_stmt_1321/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1320/do_while_stmt_1321/loop_taken/$entry
      -- 
    outputPort_4_Daemon_CP_1900_elements(5) <= outputPort_4_Daemon_CP_1900_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	158 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1320/do_while_stmt_1321/loop_body_done
      -- 
    outputPort_4_Daemon_CP_1900_elements(6) <= outputPort_4_Daemon_CP_1900_elements(158);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	38 
    -- CP-element group 7: 	59 
    -- CP-element group 7: 	80 
    -- CP-element group 7: 	101 
    -- CP-element group 7: 	122 
    -- CP-element group 7: 	141 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/back_edge_to_loop_body
      -- 
    outputPort_4_Daemon_CP_1900_elements(7) <= outputPort_4_Daemon_CP_1900_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	143 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	40 
    -- CP-element group 8: 	61 
    -- CP-element group 8: 	82 
    -- CP-element group 8: 	103 
    -- CP-element group 8: 	124 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/first_time_through_loop_body
      -- 
    outputPort_4_Daemon_CP_1900_elements(8) <= outputPort_4_Daemon_CP_1900_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	157 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	33 
    -- CP-element group 9: 	53 
    -- CP-element group 9: 	54 
    -- CP-element group 9: 	74 
    -- CP-element group 9: 	75 
    -- CP-element group 9: 	95 
    -- CP-element group 9: 	96 
    -- CP-element group 9: 	116 
    -- CP-element group 9: 	117 
    -- CP-element group 9: 	135 
    -- CP-element group 9: 	136 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/$entry
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	157 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/condition_evaluated
      -- 
    condition_evaluated_1924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(10), ack => do_while_stmt_1321_branch_req_0); -- 
    outputPort_4_Daemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(157) & outputPort_4_Daemon_CP_1900_elements(14);
      gj_outputPort_4_Daemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	32 
    -- CP-element group 11: 	53 
    -- CP-element group 11: 	74 
    -- CP-element group 11: 	95 
    -- CP-element group 11: 	116 
    -- CP-element group 11: 	135 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	55 
    -- CP-element group 11: 	76 
    -- CP-element group 11: 	97 
    -- CP-element group 11: 	118 
    -- CP-element group 11: 	137 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/aggregated_phi_sample_req
      -- 
    outputPort_4_Daemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(15) & outputPort_4_Daemon_CP_1900_elements(32) & outputPort_4_Daemon_CP_1900_elements(53) & outputPort_4_Daemon_CP_1900_elements(74) & outputPort_4_Daemon_CP_1900_elements(95) & outputPort_4_Daemon_CP_1900_elements(116) & outputPort_4_Daemon_CP_1900_elements(135) & outputPort_4_Daemon_CP_1900_elements(14);
      gj_outputPort_4_Daemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	56 
    -- CP-element group 12: 	77 
    -- CP-element group 12: 	98 
    -- CP-element group 12: 	119 
    -- CP-element group 12: 	138 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	158 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	32 
    -- CP-element group 12: 	53 
    -- CP-element group 12: 	74 
    -- CP-element group 12: 	95 
    -- CP-element group 12: 	116 
    -- CP-element group 12: 	135 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1337_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1327_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1332_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1342_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1347_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1351_sample_completed_
      -- 
    outputPort_4_Daemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(17) & outputPort_4_Daemon_CP_1900_elements(35) & outputPort_4_Daemon_CP_1900_elements(56) & outputPort_4_Daemon_CP_1900_elements(77) & outputPort_4_Daemon_CP_1900_elements(98) & outputPort_4_Daemon_CP_1900_elements(119) & outputPort_4_Daemon_CP_1900_elements(138);
      gj_outputPort_4_Daemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	33 
    -- CP-element group 13: 	54 
    -- CP-element group 13: 	75 
    -- CP-element group 13: 	96 
    -- CP-element group 13: 	117 
    -- CP-element group 13: 	136 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	36 
    -- CP-element group 13: 	57 
    -- CP-element group 13: 	78 
    -- CP-element group 13: 	99 
    -- CP-element group 13: 	120 
    -- CP-element group 13: 	139 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_update_start__ps
      -- 
    outputPort_4_Daemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(16) & outputPort_4_Daemon_CP_1900_elements(33) & outputPort_4_Daemon_CP_1900_elements(54) & outputPort_4_Daemon_CP_1900_elements(75) & outputPort_4_Daemon_CP_1900_elements(96) & outputPort_4_Daemon_CP_1900_elements(117) & outputPort_4_Daemon_CP_1900_elements(136);
      gj_outputPort_4_Daemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	37 
    -- CP-element group 14: 	58 
    -- CP-element group 14: 	79 
    -- CP-element group 14: 	100 
    -- CP-element group 14: 	121 
    -- CP-element group 14: 	140 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/aggregated_phi_update_ack
      -- 
    outputPort_4_Daemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(18) & outputPort_4_Daemon_CP_1900_elements(37) & outputPort_4_Daemon_CP_1900_elements(58) & outputPort_4_Daemon_CP_1900_elements(79) & outputPort_4_Daemon_CP_1900_elements(100) & outputPort_4_Daemon_CP_1900_elements(121) & outputPort_4_Daemon_CP_1900_elements(140);
      gj_outputPort_4_Daemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	155 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(155);
      gj_outputPort_4_Daemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	154 
    -- CP-element group 18: 	14 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_update_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(19) <= outputPort_4_Daemon_CP_1900_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_loopback_sample_req_ps
      -- CP-element group 20: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_loopback_sample_req
      -- 
    phi_stmt_1323_loopback_sample_req_1939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1323_loopback_sample_req_1939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(20), ack => phi_stmt_1323_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_entry_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(21) <= outputPort_4_Daemon_CP_1900_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_entry_sample_req_ps
      -- CP-element group 22: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_entry_sample_req
      -- 
    phi_stmt_1323_entry_sample_req_1942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1323_entry_sample_req_1942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(22), ack => phi_stmt_1323_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_phi_mux_ack_ps
      -- CP-element group 23: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_phi_mux_ack
      -- 
    phi_stmt_1323_phi_mux_ack_1945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1323_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_8_1325_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_8_1325_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_8_1325_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_8_1325_sample_start_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_8_1325_update_start_
      -- CP-element group 25: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_8_1325_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_8_1325_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(26) <= outputPort_4_Daemon_CP_1900_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_8_1325_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_1900_elements(25), ack => outputPort_4_Daemon_CP_1900_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_down_counter_1326_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_down_counter_1326_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_down_counter_1326_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_down_counter_1326_Sample/req
      -- 
    req_1966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(28), ack => next_down_counter_1438_1326_buf_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_down_counter_1326_update_start_
      -- CP-element group 29: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_down_counter_1326_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_down_counter_1326_Update/req
      -- CP-element group 29: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_down_counter_1326_Update/$entry
      -- 
    req_1971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(29), ack => next_down_counter_1438_1326_buf_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_down_counter_1326_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_down_counter_1326_Sample/ack
      -- CP-element group 30: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_down_counter_1326_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_down_counter_1326_Sample/$exit
      -- 
    ack_1967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_1438_1326_buf_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_down_counter_1326_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_down_counter_1326_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_down_counter_1326_Update/ack
      -- CP-element group 31: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_down_counter_1326_Update/$exit
      -- 
    ack_1972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_down_counter_1438_1326_buf_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	12 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	11 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1327_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	9 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	155 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	13 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1327_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(155);
      gj_outputPort_4_Daemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	11 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1327_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(34) <= outputPort_4_Daemon_CP_1900_elements(11);
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1327_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(35) is bound as output of CP function.
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	13 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1327_update_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(36) <= outputPort_4_Daemon_CP_1900_elements(13);
    -- CP-element group 37:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	154 
    -- CP-element group 37: 	14 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1327_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1327_update_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	7 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1327_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(38) <= outputPort_4_Daemon_CP_1900_elements(7);
    -- CP-element group 39:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1327_loopback_sample_req_ps
      -- CP-element group 39: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1327_loopback_sample_req
      -- 
    phi_stmt_1327_loopback_sample_req_1983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1327_loopback_sample_req_1983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(39), ack => phi_stmt_1327_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	8 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1327_entry_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(40) <= outputPort_4_Daemon_CP_1900_elements(8);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1327_entry_sample_req
      -- CP-element group 41: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1327_entry_sample_req_ps
      -- 
    phi_stmt_1327_entry_sample_req_1986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1327_entry_sample_req_1986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(41), ack => phi_stmt_1327_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(41) is bound as output of CP function.
    -- CP-element group 42:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1327_phi_mux_ack_ps
      -- CP-element group 42: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1327_phi_mux_ack
      -- 
    phi_stmt_1327_phi_mux_ack_1989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1327_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (4) 
      -- CP-element group 43: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1329_sample_start__ps
      -- CP-element group 43: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1329_sample_completed__ps
      -- CP-element group 43: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1329_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1329_sample_start_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1329_update_start_
      -- CP-element group 44: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1329_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(44) is bound as output of CP function.
    -- CP-element group 45:  join  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1329_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(45) <= outputPort_4_Daemon_CP_1900_elements(46);
    -- CP-element group 46:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	45 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1329_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(46) is a control-delay.
    cp_element_46_delay: control_delay_element  generic map(name => " 46_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_1900_elements(44), ack => outputPort_4_Daemon_CP_1900_elements(46), clk => clk, reset =>reset);
    -- CP-element group 47:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_1_4_1331_sample_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_1_4_1331_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: marked-predecessors 
    -- CP-element group 49: 	52 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_1_4_1331_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_1_4_1331_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_1_4_1331_Sample/rr
      -- 
    rr_2010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(49), ack => RPIPE_noblock_obuf_1_4_1331_inst_req_0); -- 
    outputPort_4_Daemon_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(47) & outputPort_4_Daemon_CP_1900_elements(52);
      gj_outputPort_4_Daemon_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: 	51 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_1_4_1331_update_start_
      -- CP-element group 50: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_1_4_1331_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_1_4_1331_Update/cr
      -- 
    cr_2015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(50), ack => RPIPE_noblock_obuf_1_4_1331_inst_req_1); -- 
    outputPort_4_Daemon_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(48) & outputPort_4_Daemon_CP_1900_elements(51);
      gj_outputPort_4_Daemon_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	50 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_1_4_1331_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_1_4_1331_sample_completed__ps
      -- CP-element group 51: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_1_4_1331_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_1_4_1331_Sample/ra
      -- 
    ra_2011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_4_1331_inst_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(51)); -- 
    -- CP-element group 52:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: marked-successors 
    -- CP-element group 52: 	49 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_1_4_1331_Update/ca
      -- CP-element group 52: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_1_4_1331_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_1_4_1331_update_completed__ps
      -- CP-element group 52: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_1_4_1331_Update/$exit
      -- 
    ca_2016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_1_4_1331_inst_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(52)); -- 
    -- CP-element group 53:  join  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	9 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	12 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	11 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1332_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	9 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	155 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	13 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1332_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(155);
      gj_outputPort_4_Daemon_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	11 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1332_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(55) <= outputPort_4_Daemon_CP_1900_elements(11);
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	12 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1332_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(56) is bound as output of CP function.
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	13 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1332_update_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(57) <= outputPort_4_Daemon_CP_1900_elements(13);
    -- CP-element group 58:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	154 
    -- CP-element group 58: 	14 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1332_update_completed__ps
      -- CP-element group 58: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1332_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	7 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1332_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(59) <= outputPort_4_Daemon_CP_1900_elements(7);
    -- CP-element group 60:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1332_loopback_sample_req_ps
      -- CP-element group 60: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1332_loopback_sample_req
      -- 
    phi_stmt_1332_loopback_sample_req_2027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1332_loopback_sample_req_2027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(60), ack => phi_stmt_1332_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	8 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1332_entry_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(61) <= outputPort_4_Daemon_CP_1900_elements(8);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1332_entry_sample_req
      -- CP-element group 62: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1332_entry_sample_req_ps
      -- 
    phi_stmt_1332_entry_sample_req_2030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1332_entry_sample_req_2030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(62), ack => phi_stmt_1332_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1332_phi_mux_ack_ps
      -- CP-element group 63: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1332_phi_mux_ack
      -- 
    phi_stmt_1332_phi_mux_ack_2033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1332_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(63)); -- 
    -- CP-element group 64:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (4) 
      -- CP-element group 64: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1334_sample_completed__ps
      -- CP-element group 64: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1334_sample_start__ps
      -- CP-element group 64: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1334_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1334_sample_start_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1334_update_start__ps
      -- CP-element group 65: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1334_update_start_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(65) is bound as output of CP function.
    -- CP-element group 66:  join  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1334_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(66) <= outputPort_4_Daemon_CP_1900_elements(67);
    -- CP-element group 67:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	66 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1334_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(67) is a control-delay.
    cp_element_67_delay: control_delay_element  generic map(name => " 67_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_1900_elements(65), ack => outputPort_4_Daemon_CP_1900_elements(67), clk => clk, reset =>reset);
    -- CP-element group 68:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_2_4_1336_sample_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_2_4_1336_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(69) is bound as output of CP function.
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	73 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_2_4_1336_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_2_4_1336_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_2_4_1336_sample_start_
      -- 
    rr_2054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(70), ack => RPIPE_noblock_obuf_2_4_1336_inst_req_0); -- 
    outputPort_4_Daemon_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(68) & outputPort_4_Daemon_CP_1900_elements(73);
      gj_outputPort_4_Daemon_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: 	72 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_2_4_1336_Update/cr
      -- CP-element group 71: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_2_4_1336_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_2_4_1336_update_start_
      -- 
    cr_2059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(71), ack => RPIPE_noblock_obuf_2_4_1336_inst_req_1); -- 
    outputPort_4_Daemon_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(69) & outputPort_4_Daemon_CP_1900_elements(72);
      gj_outputPort_4_Daemon_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	71 
    -- CP-element group 72:  members (4) 
      -- CP-element group 72: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_2_4_1336_Sample/ra
      -- CP-element group 72: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_2_4_1336_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_2_4_1336_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_2_4_1336_sample_completed__ps
      -- 
    ra_2055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_4_1336_inst_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(72)); -- 
    -- CP-element group 73:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: marked-successors 
    -- CP-element group 73: 	70 
    -- CP-element group 73:  members (4) 
      -- CP-element group 73: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_2_4_1336_Update/ca
      -- CP-element group 73: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_2_4_1336_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_2_4_1336_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_2_4_1336_update_completed__ps
      -- 
    ca_2060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_2_4_1336_inst_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(73)); -- 
    -- CP-element group 74:  join  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	9 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	12 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	11 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1337_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	9 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	155 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	13 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1337_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(155);
      gj_outputPort_4_Daemon_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	11 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1337_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(76) <= outputPort_4_Daemon_CP_1900_elements(11);
    -- CP-element group 77:  join  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	12 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1337_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(77) is bound as output of CP function.
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	13 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1337_update_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(78) <= outputPort_4_Daemon_CP_1900_elements(13);
    -- CP-element group 79:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	154 
    -- CP-element group 79: 	14 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1337_update_completed__ps
      -- CP-element group 79: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1337_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	7 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1337_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(80) <= outputPort_4_Daemon_CP_1900_elements(7);
    -- CP-element group 81:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1337_loopback_sample_req
      -- CP-element group 81: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1337_loopback_sample_req_ps
      -- 
    phi_stmt_1337_loopback_sample_req_2071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1337_loopback_sample_req_2071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(81), ack => phi_stmt_1337_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	8 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1337_entry_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(82) <= outputPort_4_Daemon_CP_1900_elements(8);
    -- CP-element group 83:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1337_entry_sample_req
      -- CP-element group 83: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1337_entry_sample_req_ps
      -- 
    phi_stmt_1337_entry_sample_req_2074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1337_entry_sample_req_2074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(83), ack => phi_stmt_1337_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(83) is bound as output of CP function.
    -- CP-element group 84:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1337_phi_mux_ack_ps
      -- CP-element group 84: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1337_phi_mux_ack
      -- 
    phi_stmt_1337_phi_mux_ack_2077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1337_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(84)); -- 
    -- CP-element group 85:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (4) 
      -- CP-element group 85: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1339_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1339_sample_completed__ps
      -- CP-element group 85: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1339_sample_start__ps
      -- CP-element group 85: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1339_sample_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1339_update_start__ps
      -- CP-element group 86: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1339_update_start_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(86) is bound as output of CP function.
    -- CP-element group 87:  join  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1339_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(87) <= outputPort_4_Daemon_CP_1900_elements(88);
    -- CP-element group 88:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	87 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1339_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(88) is a control-delay.
    cp_element_88_delay: control_delay_element  generic map(name => " 88_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_1900_elements(86), ack => outputPort_4_Daemon_CP_1900_elements(88), clk => clk, reset =>reset);
    -- CP-element group 89:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_3_4_1341_sample_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(89) is bound as output of CP function.
    -- CP-element group 90:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_3_4_1341_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(90) is bound as output of CP function.
    -- CP-element group 91:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: marked-predecessors 
    -- CP-element group 91: 	94 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_3_4_1341_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_3_4_1341_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_3_4_1341_Sample/$entry
      -- 
    rr_2098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(91), ack => RPIPE_noblock_obuf_3_4_1341_inst_req_0); -- 
    outputPort_4_Daemon_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(89) & outputPort_4_Daemon_CP_1900_elements(94);
      gj_outputPort_4_Daemon_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	93 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_3_4_1341_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_3_4_1341_update_start_
      -- CP-element group 92: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_3_4_1341_Update/$entry
      -- 
    cr_2103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(92), ack => RPIPE_noblock_obuf_3_4_1341_inst_req_1); -- 
    outputPort_4_Daemon_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(90) & outputPort_4_Daemon_CP_1900_elements(93);
      gj_outputPort_4_Daemon_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	92 
    -- CP-element group 93:  members (4) 
      -- CP-element group 93: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_3_4_1341_sample_completed__ps
      -- CP-element group 93: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_3_4_1341_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_3_4_1341_Sample/ra
      -- CP-element group 93: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_3_4_1341_Sample/$exit
      -- 
    ra_2099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_4_1341_inst_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(93)); -- 
    -- CP-element group 94:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: successors 
    -- CP-element group 94: marked-successors 
    -- CP-element group 94: 	91 
    -- CP-element group 94:  members (4) 
      -- CP-element group 94: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_3_4_1341_update_completed__ps
      -- CP-element group 94: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_3_4_1341_Update/ca
      -- CP-element group 94: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_3_4_1341_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_3_4_1341_Update/$exit
      -- 
    ca_2104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_3_4_1341_inst_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(94)); -- 
    -- CP-element group 95:  join  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	9 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	12 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	11 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1342_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	9 
    -- CP-element group 96: marked-predecessors 
    -- CP-element group 96: 	155 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	13 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1342_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "outputPort_4_Daemon_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(155);
      gj_outputPort_4_Daemon_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	11 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1342_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(97) <= outputPort_4_Daemon_CP_1900_elements(11);
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	12 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1342_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(98) is bound as output of CP function.
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	13 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1342_update_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(99) <= outputPort_4_Daemon_CP_1900_elements(13);
    -- CP-element group 100:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	154 
    -- CP-element group 100: 	14 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1342_update_completed__ps
      -- CP-element group 100: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1342_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(100) is bound as output of CP function.
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	7 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1342_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(101) <= outputPort_4_Daemon_CP_1900_elements(7);
    -- CP-element group 102:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1342_loopback_sample_req_ps
      -- CP-element group 102: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1342_loopback_sample_req
      -- 
    phi_stmt_1342_loopback_sample_req_2115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1342_loopback_sample_req_2115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(102), ack => phi_stmt_1342_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(102) is bound as output of CP function.
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	8 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1342_entry_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(103) <= outputPort_4_Daemon_CP_1900_elements(8);
    -- CP-element group 104:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1342_entry_sample_req_ps
      -- CP-element group 104: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1342_entry_sample_req
      -- 
    phi_stmt_1342_entry_sample_req_2118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1342_entry_sample_req_2118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(104), ack => phi_stmt_1342_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(104) is bound as output of CP function.
    -- CP-element group 105:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1342_phi_mux_ack_ps
      -- CP-element group 105: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1342_phi_mux_ack
      -- 
    phi_stmt_1342_phi_mux_ack_2121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1342_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(105)); -- 
    -- CP-element group 106:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (4) 
      -- CP-element group 106: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1344_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1344_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1344_sample_completed__ps
      -- CP-element group 106: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1344_sample_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1344_update_start_
      -- CP-element group 107: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1344_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(107) is bound as output of CP function.
    -- CP-element group 108:  join  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	109 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1344_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(108) <= outputPort_4_Daemon_CP_1900_elements(109);
    -- CP-element group 109:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	108 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_33_1344_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(109) is a control-delay.
    cp_element_109_delay: control_delay_element  generic map(name => " 109_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_1900_elements(107), ack => outputPort_4_Daemon_CP_1900_elements(109), clk => clk, reset =>reset);
    -- CP-element group 110:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_4_4_1346_sample_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(110) is bound as output of CP function.
    -- CP-element group 111:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_4_4_1346_update_start__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(111) is bound as output of CP function.
    -- CP-element group 112:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	115 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_4_4_1346_Sample/rr
      -- CP-element group 112: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_4_4_1346_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_4_4_1346_sample_start_
      -- 
    rr_2142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(112), ack => RPIPE_noblock_obuf_4_4_1346_inst_req_0); -- 
    outputPort_4_Daemon_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(110) & outputPort_4_Daemon_CP_1900_elements(115);
      gj_outputPort_4_Daemon_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: 	114 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_4_4_1346_Update/cr
      -- CP-element group 113: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_4_4_1346_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_4_4_1346_update_start_
      -- 
    cr_2147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(113), ack => RPIPE_noblock_obuf_4_4_1346_inst_req_1); -- 
    outputPort_4_Daemon_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(111) & outputPort_4_Daemon_CP_1900_elements(114);
      gj_outputPort_4_Daemon_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	113 
    -- CP-element group 114:  members (4) 
      -- CP-element group 114: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_4_4_1346_Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_4_4_1346_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_4_4_1346_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_4_4_1346_sample_completed__ps
      -- 
    ra_2143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_4_1346_inst_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(114)); -- 
    -- CP-element group 115:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	112 
    -- CP-element group 115:  members (4) 
      -- CP-element group 115: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_4_4_1346_Update/ca
      -- CP-element group 115: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_4_4_1346_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_4_4_1346_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_noblock_obuf_4_4_1346_update_completed__ps
      -- 
    ca_2148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_noblock_obuf_4_4_1346_inst_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(115)); -- 
    -- CP-element group 116:  join  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	9 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	12 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	11 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1347_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  transition  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	9 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	155 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	13 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1347_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(155);
      gj_outputPort_4_Daemon_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	11 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1347_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(118) <= outputPort_4_Daemon_CP_1900_elements(11);
    -- CP-element group 119:  join  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	12 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1347_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(119) is bound as output of CP function.
    -- CP-element group 120:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	13 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1347_update_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(120) <= outputPort_4_Daemon_CP_1900_elements(13);
    -- CP-element group 121:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	154 
    -- CP-element group 121: 	14 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1347_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1347_update_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(121) is bound as output of CP function.
    -- CP-element group 122:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	7 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1347_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(122) <= outputPort_4_Daemon_CP_1900_elements(7);
    -- CP-element group 123:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1347_loopback_sample_req
      -- CP-element group 123: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1347_loopback_sample_req_ps
      -- 
    phi_stmt_1347_loopback_sample_req_2159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1347_loopback_sample_req_2159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(123), ack => phi_stmt_1347_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(123) is bound as output of CP function.
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	8 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1347_entry_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(124) <= outputPort_4_Daemon_CP_1900_elements(8);
    -- CP-element group 125:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1347_entry_sample_req
      -- CP-element group 125: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1347_entry_sample_req_ps
      -- 
    phi_stmt_1347_entry_sample_req_2162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1347_entry_sample_req_2162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(125), ack => phi_stmt_1347_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(125) is bound as output of CP function.
    -- CP-element group 126:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1347_phi_mux_ack
      -- CP-element group 126: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1347_phi_mux_ack_ps
      -- 
    phi_stmt_1347_phi_mux_ack_2165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1347_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(126)); -- 
    -- CP-element group 127:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (4) 
      -- CP-element group 127: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_3_1349_sample_start__ps
      -- CP-element group 127: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_3_1349_sample_completed__ps
      -- CP-element group 127: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_3_1349_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_3_1349_sample_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(127) is bound as output of CP function.
    -- CP-element group 128:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_3_1349_update_start__ps
      -- CP-element group 128: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_3_1349_update_start_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(128) is bound as output of CP function.
    -- CP-element group 129:  join  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	130 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_3_1349_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(129) <= outputPort_4_Daemon_CP_1900_elements(130);
    -- CP-element group 130:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	129 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_3_1349_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(130) is a control-delay.
    cp_element_130_delay: control_delay_element  generic map(name => " 130_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_1900_elements(128), ack => outputPort_4_Daemon_CP_1900_elements(130), clk => clk, reset =>reset);
    -- CP-element group 131:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (4) 
      -- CP-element group 131: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_active_packet_1350_sample_start__ps
      -- CP-element group 131: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_active_packet_1350_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_active_packet_1350_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_active_packet_1350_Sample/req
      -- 
    req_2186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(131), ack => next_active_packet_1414_1350_buf_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(131) is bound as output of CP function.
    -- CP-element group 132:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (4) 
      -- CP-element group 132: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_active_packet_1350_update_start__ps
      -- CP-element group 132: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_active_packet_1350_update_start_
      -- CP-element group 132: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_active_packet_1350_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_active_packet_1350_Update/req
      -- 
    req_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(132), ack => next_active_packet_1414_1350_buf_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(132) is bound as output of CP function.
    -- CP-element group 133:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_active_packet_1350_sample_completed__ps
      -- CP-element group 133: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_active_packet_1350_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_active_packet_1350_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_active_packet_1350_Sample/ack
      -- 
    ack_2187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_1414_1350_buf_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(133)); -- 
    -- CP-element group 134:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_active_packet_1350_update_completed__ps
      -- CP-element group 134: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_active_packet_1350_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_active_packet_1350_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_active_packet_1350_Update/ack
      -- 
    ack_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_active_packet_1414_1350_buf_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(134)); -- 
    -- CP-element group 135:  join  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	9 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	12 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	11 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1351_sample_start_
      -- 
    outputPort_4_Daemon_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	9 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	155 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	13 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1351_update_start_
      -- 
    outputPort_4_Daemon_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(9) & outputPort_4_Daemon_CP_1900_elements(155);
      gj_outputPort_4_Daemon_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	11 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1351_sample_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(137) <= outputPort_4_Daemon_CP_1900_elements(11);
    -- CP-element group 138:  join  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	12 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1351_sample_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(138) is bound as output of CP function.
    -- CP-element group 139:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	13 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1351_update_start__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(139) <= outputPort_4_Daemon_CP_1900_elements(13);
    -- CP-element group 140:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	154 
    -- CP-element group 140: 	14 
    -- CP-element group 140:  members (2) 
      -- CP-element group 140: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1351_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1351_update_completed__ps
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(140) is bound as output of CP function.
    -- CP-element group 141:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	7 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1351_loopback_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(141) <= outputPort_4_Daemon_CP_1900_elements(7);
    -- CP-element group 142:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1351_loopback_sample_req
      -- CP-element group 142: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1351_loopback_sample_req_ps
      -- 
    phi_stmt_1351_loopback_sample_req_2203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1351_loopback_sample_req_2203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(142), ack => phi_stmt_1351_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(142) is bound as output of CP function.
    -- CP-element group 143:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	8 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1351_entry_trigger
      -- 
    outputPort_4_Daemon_CP_1900_elements(143) <= outputPort_4_Daemon_CP_1900_elements(8);
    -- CP-element group 144:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1351_entry_sample_req
      -- CP-element group 144: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1351_entry_sample_req_ps
      -- 
    phi_stmt_1351_entry_sample_req_2206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1351_entry_sample_req_2206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(144), ack => phi_stmt_1351_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1351_phi_mux_ack
      -- CP-element group 145: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1351_phi_mux_ack_ps
      -- 
    phi_stmt_1351_phi_mux_ack_2209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1351_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(145)); -- 
    -- CP-element group 146:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (4) 
      -- CP-element group 146: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_3_1353_sample_start__ps
      -- CP-element group 146: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_3_1353_sample_completed__ps
      -- CP-element group 146: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_3_1353_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_3_1353_sample_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(146) is bound as output of CP function.
    -- CP-element group 147:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (2) 
      -- CP-element group 147: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_3_1353_update_start__ps
      -- CP-element group 147: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_3_1353_update_start_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(147) is bound as output of CP function.
    -- CP-element group 148:  join  transition  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	149 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (1) 
      -- CP-element group 148: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_3_1353_update_completed__ps
      -- 
    outputPort_4_Daemon_CP_1900_elements(148) <= outputPort_4_Daemon_CP_1900_elements(149);
    -- CP-element group 149:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	148 
    -- CP-element group 149:  members (1) 
      -- CP-element group 149: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_ZERO_3_1353_update_completed_
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(149) is a control-delay.
    cp_element_149_delay: control_delay_element  generic map(name => " 149_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_1900_elements(147), ack => outputPort_4_Daemon_CP_1900_elements(149), clk => clk, reset =>reset);
    -- CP-element group 150:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (4) 
      -- CP-element group 150: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_pkt_priority_1354_sample_start__ps
      -- CP-element group 150: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_pkt_priority_1354_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_pkt_priority_1354_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_pkt_priority_1354_Sample/req
      -- 
    req_2230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(150), ack => next_pkt_priority_1414_1354_buf_req_0); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(150) is bound as output of CP function.
    -- CP-element group 151:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (4) 
      -- CP-element group 151: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_pkt_priority_1354_update_start__ps
      -- CP-element group 151: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_pkt_priority_1354_update_start_
      -- CP-element group 151: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_pkt_priority_1354_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_pkt_priority_1354_Update/req
      -- 
    req_2235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(151), ack => next_pkt_priority_1414_1354_buf_req_1); -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(151) is bound as output of CP function.
    -- CP-element group 152:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (4) 
      -- CP-element group 152: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_pkt_priority_1354_sample_completed__ps
      -- CP-element group 152: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_pkt_priority_1354_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_pkt_priority_1354_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_pkt_priority_1354_Sample/ack
      -- 
    ack_2231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pkt_priority_1414_1354_buf_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(152)); -- 
    -- CP-element group 153:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (4) 
      -- CP-element group 153: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_pkt_priority_1354_update_completed__ps
      -- CP-element group 153: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_pkt_priority_1354_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_pkt_priority_1354_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_next_pkt_priority_1354_Update/ack
      -- 
    ack_2236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_pkt_priority_1414_1354_buf_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	18 
    -- CP-element group 154: 	37 
    -- CP-element group 154: 	58 
    -- CP-element group 154: 	79 
    -- CP-element group 154: 	100 
    -- CP-element group 154: 	121 
    -- CP-element group 154: 	140 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/WPIPE_out_data_4_1534_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/WPIPE_out_data_4_1534_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/WPIPE_out_data_4_1534_Sample/req
      -- 
    req_2245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(154), ack => WPIPE_out_data_4_1534_inst_req_0); -- 
    outputPort_4_Daemon_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 7,1 => 7,2 => 7,3 => 7,4 => 7,5 => 7,6 => 7,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(18) & outputPort_4_Daemon_CP_1900_elements(37) & outputPort_4_Daemon_CP_1900_elements(58) & outputPort_4_Daemon_CP_1900_elements(79) & outputPort_4_Daemon_CP_1900_elements(100) & outputPort_4_Daemon_CP_1900_elements(121) & outputPort_4_Daemon_CP_1900_elements(140) & outputPort_4_Daemon_CP_1900_elements(156);
      gj_outputPort_4_Daemon_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	16 
    -- CP-element group 155: 	33 
    -- CP-element group 155: 	54 
    -- CP-element group 155: 	75 
    -- CP-element group 155: 	96 
    -- CP-element group 155: 	117 
    -- CP-element group 155: 	136 
    -- CP-element group 155:  members (6) 
      -- CP-element group 155: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/WPIPE_out_data_4_1534_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/WPIPE_out_data_4_1534_update_start_
      -- CP-element group 155: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/WPIPE_out_data_4_1534_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/WPIPE_out_data_4_1534_Sample/ack
      -- CP-element group 155: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/WPIPE_out_data_4_1534_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/WPIPE_out_data_4_1534_Update/req
      -- 
    ack_2246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_4_1534_inst_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(155)); -- 
    req_2250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => outputPort_4_Daemon_CP_1900_elements(155), ack => WPIPE_out_data_4_1534_inst_req_1); -- 
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	154 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/WPIPE_out_data_4_1534_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/WPIPE_out_data_4_1534_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/WPIPE_out_data_4_1534_Update/ack
      -- 
    ack_2251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_out_data_4_1534_inst_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(156)); -- 
    -- CP-element group 157:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	9 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	10 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group outputPort_4_Daemon_CP_1900_elements(157) is a control-delay.
    cp_element_157_delay: control_delay_element  generic map(name => " 157_delay", delay_value => 1)  port map(req => outputPort_4_Daemon_CP_1900_elements(9), ack => outputPort_4_Daemon_CP_1900_elements(157), clk => clk, reset =>reset);
    -- CP-element group 158:  join  transition  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: 	12 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	6 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/$exit
      -- 
    outputPort_4_Daemon_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "outputPort_4_Daemon_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= outputPort_4_Daemon_CP_1900_elements(156) & outputPort_4_Daemon_CP_1900_elements(12);
      gj_outputPort_4_Daemon_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	5 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (2) 
      -- CP-element group 159: 	 branch_block_stmt_1320/do_while_stmt_1321/loop_exit/$exit
      -- CP-element group 159: 	 branch_block_stmt_1320/do_while_stmt_1321/loop_exit/ack
      -- 
    ack_2256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1321_branch_ack_0, ack => outputPort_4_Daemon_CP_1900_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	5 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (2) 
      -- CP-element group 160: 	 branch_block_stmt_1320/do_while_stmt_1321/loop_taken/$exit
      -- CP-element group 160: 	 branch_block_stmt_1320/do_while_stmt_1321/loop_taken/ack
      -- 
    ack_2260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1321_branch_ack_1, ack => outputPort_4_Daemon_CP_1900_elements(160)); -- 
    -- CP-element group 161:  transition  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	3 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	1 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_1320/do_while_stmt_1321/$exit
      -- 
    outputPort_4_Daemon_CP_1900_elements(161) <= outputPort_4_Daemon_CP_1900_elements(3);
    outputPort_4_Daemon_do_while_stmt_1321_terminator_2261: loop_terminator -- 
      generic map (name => " outputPort_4_Daemon_do_while_stmt_1321_terminator_2261", max_iterations_in_flight =>7) 
      port map(loop_body_exit => outputPort_4_Daemon_CP_1900_elements(6),loop_continue => outputPort_4_Daemon_CP_1900_elements(160),loop_terminate => outputPort_4_Daemon_CP_1900_elements(159),loop_back => outputPort_4_Daemon_CP_1900_elements(4),loop_exit => outputPort_4_Daemon_CP_1900_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1323_phi_seq_1973_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_1900_elements(21);
      outputPort_4_Daemon_CP_1900_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(24);
      outputPort_4_Daemon_CP_1900_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(26);
      outputPort_4_Daemon_CP_1900_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_1900_elements(19);
      outputPort_4_Daemon_CP_1900_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(30);
      outputPort_4_Daemon_CP_1900_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(31);
      outputPort_4_Daemon_CP_1900_elements(20) <= phi_mux_reqs(1);
      phi_stmt_1323_phi_seq_1973 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1323_phi_seq_1973") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_1900_elements(11), 
          phi_sample_ack => outputPort_4_Daemon_CP_1900_elements(17), 
          phi_update_req => outputPort_4_Daemon_CP_1900_elements(13), 
          phi_update_ack => outputPort_4_Daemon_CP_1900_elements(18), 
          phi_mux_ack => outputPort_4_Daemon_CP_1900_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1327_phi_seq_2017_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_1900_elements(40);
      outputPort_4_Daemon_CP_1900_elements(43)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(43);
      outputPort_4_Daemon_CP_1900_elements(44)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(45);
      outputPort_4_Daemon_CP_1900_elements(41) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_1900_elements(38);
      outputPort_4_Daemon_CP_1900_elements(47)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(51);
      outputPort_4_Daemon_CP_1900_elements(48)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(52);
      outputPort_4_Daemon_CP_1900_elements(39) <= phi_mux_reqs(1);
      phi_stmt_1327_phi_seq_2017 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1327_phi_seq_2017") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_1900_elements(34), 
          phi_sample_ack => outputPort_4_Daemon_CP_1900_elements(35), 
          phi_update_req => outputPort_4_Daemon_CP_1900_elements(36), 
          phi_update_ack => outputPort_4_Daemon_CP_1900_elements(37), 
          phi_mux_ack => outputPort_4_Daemon_CP_1900_elements(42), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1332_phi_seq_2061_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_1900_elements(61);
      outputPort_4_Daemon_CP_1900_elements(64)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(64);
      outputPort_4_Daemon_CP_1900_elements(65)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(66);
      outputPort_4_Daemon_CP_1900_elements(62) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_1900_elements(59);
      outputPort_4_Daemon_CP_1900_elements(68)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(72);
      outputPort_4_Daemon_CP_1900_elements(69)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(73);
      outputPort_4_Daemon_CP_1900_elements(60) <= phi_mux_reqs(1);
      phi_stmt_1332_phi_seq_2061 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1332_phi_seq_2061") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_1900_elements(55), 
          phi_sample_ack => outputPort_4_Daemon_CP_1900_elements(56), 
          phi_update_req => outputPort_4_Daemon_CP_1900_elements(57), 
          phi_update_ack => outputPort_4_Daemon_CP_1900_elements(58), 
          phi_mux_ack => outputPort_4_Daemon_CP_1900_elements(63), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1337_phi_seq_2105_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_1900_elements(82);
      outputPort_4_Daemon_CP_1900_elements(85)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(85);
      outputPort_4_Daemon_CP_1900_elements(86)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(87);
      outputPort_4_Daemon_CP_1900_elements(83) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_1900_elements(80);
      outputPort_4_Daemon_CP_1900_elements(89)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(93);
      outputPort_4_Daemon_CP_1900_elements(90)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(94);
      outputPort_4_Daemon_CP_1900_elements(81) <= phi_mux_reqs(1);
      phi_stmt_1337_phi_seq_2105 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1337_phi_seq_2105") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_1900_elements(76), 
          phi_sample_ack => outputPort_4_Daemon_CP_1900_elements(77), 
          phi_update_req => outputPort_4_Daemon_CP_1900_elements(78), 
          phi_update_ack => outputPort_4_Daemon_CP_1900_elements(79), 
          phi_mux_ack => outputPort_4_Daemon_CP_1900_elements(84), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1342_phi_seq_2149_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_1900_elements(103);
      outputPort_4_Daemon_CP_1900_elements(106)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(106);
      outputPort_4_Daemon_CP_1900_elements(107)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(108);
      outputPort_4_Daemon_CP_1900_elements(104) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_1900_elements(101);
      outputPort_4_Daemon_CP_1900_elements(110)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(114);
      outputPort_4_Daemon_CP_1900_elements(111)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(115);
      outputPort_4_Daemon_CP_1900_elements(102) <= phi_mux_reqs(1);
      phi_stmt_1342_phi_seq_2149 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1342_phi_seq_2149") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_1900_elements(97), 
          phi_sample_ack => outputPort_4_Daemon_CP_1900_elements(98), 
          phi_update_req => outputPort_4_Daemon_CP_1900_elements(99), 
          phi_update_ack => outputPort_4_Daemon_CP_1900_elements(100), 
          phi_mux_ack => outputPort_4_Daemon_CP_1900_elements(105), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1347_phi_seq_2193_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_1900_elements(124);
      outputPort_4_Daemon_CP_1900_elements(127)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(127);
      outputPort_4_Daemon_CP_1900_elements(128)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(129);
      outputPort_4_Daemon_CP_1900_elements(125) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_1900_elements(122);
      outputPort_4_Daemon_CP_1900_elements(131)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(133);
      outputPort_4_Daemon_CP_1900_elements(132)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(134);
      outputPort_4_Daemon_CP_1900_elements(123) <= phi_mux_reqs(1);
      phi_stmt_1347_phi_seq_2193 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1347_phi_seq_2193") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_1900_elements(118), 
          phi_sample_ack => outputPort_4_Daemon_CP_1900_elements(119), 
          phi_update_req => outputPort_4_Daemon_CP_1900_elements(120), 
          phi_update_ack => outputPort_4_Daemon_CP_1900_elements(121), 
          phi_mux_ack => outputPort_4_Daemon_CP_1900_elements(126), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1351_phi_seq_2237_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= outputPort_4_Daemon_CP_1900_elements(143);
      outputPort_4_Daemon_CP_1900_elements(146)<= src_sample_reqs(0);
      src_sample_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(146);
      outputPort_4_Daemon_CP_1900_elements(147)<= src_update_reqs(0);
      src_update_acks(0)  <= outputPort_4_Daemon_CP_1900_elements(148);
      outputPort_4_Daemon_CP_1900_elements(144) <= phi_mux_reqs(0);
      triggers(1)  <= outputPort_4_Daemon_CP_1900_elements(141);
      outputPort_4_Daemon_CP_1900_elements(150)<= src_sample_reqs(1);
      src_sample_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(152);
      outputPort_4_Daemon_CP_1900_elements(151)<= src_update_reqs(1);
      src_update_acks(1)  <= outputPort_4_Daemon_CP_1900_elements(153);
      outputPort_4_Daemon_CP_1900_elements(142) <= phi_mux_reqs(1);
      phi_stmt_1351_phi_seq_2237 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1351_phi_seq_2237") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => outputPort_4_Daemon_CP_1900_elements(137), 
          phi_sample_ack => outputPort_4_Daemon_CP_1900_elements(138), 
          phi_update_req => outputPort_4_Daemon_CP_1900_elements(139), 
          phi_update_ack => outputPort_4_Daemon_CP_1900_elements(140), 
          phi_mux_ack => outputPort_4_Daemon_CP_1900_elements(145), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1925_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= outputPort_4_Daemon_CP_1900_elements(7);
        preds(1)  <= outputPort_4_Daemon_CP_1900_elements(8);
        entry_tmerge_1925 : transition_merge -- 
          generic map(name => " entry_tmerge_1925")
          port map (preds => preds, symbol_out => outputPort_4_Daemon_CP_1900_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u3_u1_1379_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1385_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1392_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1398_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1444_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1452_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1460_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1468_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1474_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1481_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1489_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1496_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1507_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1513_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1520_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1526_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_1425_wire : std_logic_vector(0 downto 0);
    signal MUX_1382_wire : std_logic_vector(0 downto 0);
    signal MUX_1388_wire : std_logic_vector(0 downto 0);
    signal MUX_1395_wire : std_logic_vector(0 downto 0);
    signal MUX_1401_wire : std_logic_vector(0 downto 0);
    signal MUX_1436_wire : std_logic_vector(7 downto 0);
    signal MUX_1478_wire : std_logic_vector(31 downto 0);
    signal MUX_1485_wire : std_logic_vector(31 downto 0);
    signal MUX_1493_wire : std_logic_vector(31 downto 0);
    signal MUX_1500_wire : std_logic_vector(31 downto 0);
    signal MUX_1510_wire : std_logic_vector(0 downto 0);
    signal MUX_1516_wire : std_logic_vector(0 downto 0);
    signal MUX_1523_wire : std_logic_vector(0 downto 0);
    signal MUX_1529_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1441_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1449_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1457_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1465_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1389_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1402_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1418_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1421_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1422_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1517_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1530_wire : std_logic_vector(0 downto 0);
    signal OR_u32_u32_1486_wire : std_logic_vector(31 downto 0);
    signal OR_u32_u32_1501_wire : std_logic_vector(31 downto 0);
    signal RPIPE_noblock_obuf_1_4_1331_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_2_4_1336_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_3_4_1341_wire : std_logic_vector(32 downto 0);
    signal RPIPE_noblock_obuf_4_4_1346_wire : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1329_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1334_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1339_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_33_1344_wire_constant : std_logic_vector(32 downto 0);
    signal R_ZERO_3_1349_wire_constant : std_logic_vector(2 downto 0);
    signal R_ZERO_3_1353_wire_constant : std_logic_vector(2 downto 0);
    signal R_ZERO_8_1325_wire_constant : std_logic_vector(7 downto 0);
    signal SUB_u8_u8_1434_wire : std_logic_vector(7 downto 0);
    signal active_packet_1347 : std_logic_vector(2 downto 0);
    signal data_to_out_1503 : std_logic_vector(31 downto 0);
    signal down_counter_1323 : std_logic_vector(7 downto 0);
    signal konst_1358_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1363_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1368_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1373_wire_constant : std_logic_vector(32 downto 0);
    signal konst_1378_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1381_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1384_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1387_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1391_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1394_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1397_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1400_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1424_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1430_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1433_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1443_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1451_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1459_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1467_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1473_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1477_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1480_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1484_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1488_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1492_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1495_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1499_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1506_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1509_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1512_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1515_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1519_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1522_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1525_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1528_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1538_wire_constant : std_logic_vector(0 downto 0);
    signal next_active_packet_1414 : std_logic_vector(2 downto 0);
    signal next_active_packet_1414_1350_buffered : std_logic_vector(2 downto 0);
    signal next_down_counter_1438 : std_logic_vector(7 downto 0);
    signal next_down_counter_1438_1326_buffered : std_logic_vector(7 downto 0);
    signal next_pkt_priority_1414 : std_logic_vector(2 downto 0);
    signal next_pkt_priority_1414_1354_buffered : std_logic_vector(2 downto 0);
    signal p1_valid_1360 : std_logic_vector(0 downto 0);
    signal p2_valid_1365 : std_logic_vector(0 downto 0);
    signal p3_valid_1370 : std_logic_vector(0 downto 0);
    signal p4_valid_1375 : std_logic_vector(0 downto 0);
    signal pkt_1_e_word_1327 : std_logic_vector(32 downto 0);
    signal pkt_2_e_word_1332 : std_logic_vector(32 downto 0);
    signal pkt_3_e_word_1337 : std_logic_vector(32 downto 0);
    signal pkt_4_e_word_1342 : std_logic_vector(32 downto 0);
    signal pkt_priority_1351 : std_logic_vector(2 downto 0);
    signal read_from_1_1446 : std_logic_vector(0 downto 0);
    signal read_from_2_1454 : std_logic_vector(0 downto 0);
    signal read_from_3_1462 : std_logic_vector(0 downto 0);
    signal read_from_4_1470 : std_logic_vector(0 downto 0);
    signal send_flag_1532 : std_logic_vector(0 downto 0);
    signal slice_1476_wire : std_logic_vector(31 downto 0);
    signal slice_1483_wire : std_logic_vector(31 downto 0);
    signal slice_1491_wire : std_logic_vector(31 downto 0);
    signal slice_1498_wire : std_logic_vector(31 downto 0);
    signal started_new_packet_1427 : std_logic_vector(0 downto 0);
    signal valid_active_pkt_word_read_1404 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_ZERO_33_1329_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1334_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1339_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_33_1344_wire_constant <= "000000000000000000000000000000000";
    R_ZERO_3_1349_wire_constant <= "000";
    R_ZERO_3_1353_wire_constant <= "000";
    R_ZERO_8_1325_wire_constant <= "00000000";
    konst_1358_wire_constant <= "000000000000000000000000000100000";
    konst_1363_wire_constant <= "000000000000000000000000000100000";
    konst_1368_wire_constant <= "000000000000000000000000000100000";
    konst_1373_wire_constant <= "000000000000000000000000000100000";
    konst_1378_wire_constant <= "001";
    konst_1381_wire_constant <= "0";
    konst_1384_wire_constant <= "010";
    konst_1387_wire_constant <= "0";
    konst_1391_wire_constant <= "011";
    konst_1394_wire_constant <= "0";
    konst_1397_wire_constant <= "100";
    konst_1400_wire_constant <= "0";
    konst_1424_wire_constant <= "00000000";
    konst_1430_wire_constant <= "00111111";
    konst_1433_wire_constant <= "00000001";
    konst_1443_wire_constant <= "001";
    konst_1451_wire_constant <= "010";
    konst_1459_wire_constant <= "011";
    konst_1467_wire_constant <= "100";
    konst_1473_wire_constant <= "001";
    konst_1477_wire_constant <= "00000000000000000000000000000000";
    konst_1480_wire_constant <= "010";
    konst_1484_wire_constant <= "00000000000000000000000000000000";
    konst_1488_wire_constant <= "011";
    konst_1492_wire_constant <= "00000000000000000000000000000000";
    konst_1495_wire_constant <= "100";
    konst_1499_wire_constant <= "00000000000000000000000000000000";
    konst_1506_wire_constant <= "001";
    konst_1509_wire_constant <= "0";
    konst_1512_wire_constant <= "010";
    konst_1515_wire_constant <= "0";
    konst_1519_wire_constant <= "011";
    konst_1522_wire_constant <= "0";
    konst_1525_wire_constant <= "100";
    konst_1528_wire_constant <= "0";
    konst_1538_wire_constant <= "1";
    phi_stmt_1323: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_8_1325_wire_constant & next_down_counter_1438_1326_buffered;
      req <= phi_stmt_1323_req_0 & phi_stmt_1323_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1323",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1323_ack_0,
          idata => idata,
          odata => down_counter_1323,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1323
    phi_stmt_1327: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1329_wire_constant & RPIPE_noblock_obuf_1_4_1331_wire;
      req <= phi_stmt_1327_req_0 & phi_stmt_1327_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1327",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1327_ack_0,
          idata => idata,
          odata => pkt_1_e_word_1327,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1327
    phi_stmt_1332: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1334_wire_constant & RPIPE_noblock_obuf_2_4_1336_wire;
      req <= phi_stmt_1332_req_0 & phi_stmt_1332_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1332",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1332_ack_0,
          idata => idata,
          odata => pkt_2_e_word_1332,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1332
    phi_stmt_1337: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1339_wire_constant & RPIPE_noblock_obuf_3_4_1341_wire;
      req <= phi_stmt_1337_req_0 & phi_stmt_1337_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1337",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1337_ack_0,
          idata => idata,
          odata => pkt_3_e_word_1337,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1337
    phi_stmt_1342: Block -- phi operator 
      signal idata: std_logic_vector(65 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_33_1344_wire_constant & RPIPE_noblock_obuf_4_4_1346_wire;
      req <= phi_stmt_1342_req_0 & phi_stmt_1342_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1342",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 33) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1342_ack_0,
          idata => idata,
          odata => pkt_4_e_word_1342,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1342
    phi_stmt_1347: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_3_1349_wire_constant & next_active_packet_1414_1350_buffered;
      req <= phi_stmt_1347_req_0 & phi_stmt_1347_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1347",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1347_ack_0,
          idata => idata,
          odata => active_packet_1347,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1347
    phi_stmt_1351: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_ZERO_3_1353_wire_constant & next_pkt_priority_1414_1354_buffered;
      req <= phi_stmt_1351_req_0 & phi_stmt_1351_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1351",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1351_ack_0,
          idata => idata,
          odata => pkt_priority_1351,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1351
    -- flow-through select operator MUX_1382_inst
    MUX_1382_wire <= p1_valid_1360 when (EQ_u3_u1_1379_wire(0) /=  '0') else konst_1381_wire_constant;
    -- flow-through select operator MUX_1388_inst
    MUX_1388_wire <= p2_valid_1365 when (EQ_u3_u1_1385_wire(0) /=  '0') else konst_1387_wire_constant;
    -- flow-through select operator MUX_1395_inst
    MUX_1395_wire <= p3_valid_1370 when (EQ_u3_u1_1392_wire(0) /=  '0') else konst_1394_wire_constant;
    -- flow-through select operator MUX_1401_inst
    MUX_1401_wire <= p4_valid_1375 when (EQ_u3_u1_1398_wire(0) /=  '0') else konst_1400_wire_constant;
    -- flow-through select operator MUX_1436_inst
    MUX_1436_wire <= SUB_u8_u8_1434_wire when (valid_active_pkt_word_read_1404(0) /=  '0') else down_counter_1323;
    -- flow-through select operator MUX_1437_inst
    next_down_counter_1438 <= konst_1430_wire_constant when (started_new_packet_1427(0) /=  '0') else MUX_1436_wire;
    -- flow-through select operator MUX_1478_inst
    MUX_1478_wire <= slice_1476_wire when (EQ_u3_u1_1474_wire(0) /=  '0') else konst_1477_wire_constant;
    -- flow-through select operator MUX_1485_inst
    MUX_1485_wire <= slice_1483_wire when (EQ_u3_u1_1481_wire(0) /=  '0') else konst_1484_wire_constant;
    -- flow-through select operator MUX_1493_inst
    MUX_1493_wire <= slice_1491_wire when (EQ_u3_u1_1489_wire(0) /=  '0') else konst_1492_wire_constant;
    -- flow-through select operator MUX_1500_inst
    MUX_1500_wire <= slice_1498_wire when (EQ_u3_u1_1496_wire(0) /=  '0') else konst_1499_wire_constant;
    -- flow-through select operator MUX_1510_inst
    MUX_1510_wire <= p1_valid_1360 when (EQ_u3_u1_1507_wire(0) /=  '0') else konst_1509_wire_constant;
    -- flow-through select operator MUX_1516_inst
    MUX_1516_wire <= p2_valid_1365 when (EQ_u3_u1_1513_wire(0) /=  '0') else konst_1515_wire_constant;
    -- flow-through select operator MUX_1523_inst
    MUX_1523_wire <= p3_valid_1370 when (EQ_u3_u1_1520_wire(0) /=  '0') else konst_1522_wire_constant;
    -- flow-through select operator MUX_1529_inst
    MUX_1529_wire <= p4_valid_1375 when (EQ_u3_u1_1526_wire(0) /=  '0') else konst_1528_wire_constant;
    -- flow-through slice operator slice_1476_inst
    slice_1476_wire <= pkt_1_e_word_1327(31 downto 0);
    -- flow-through slice operator slice_1483_inst
    slice_1483_wire <= pkt_2_e_word_1332(31 downto 0);
    -- flow-through slice operator slice_1491_inst
    slice_1491_wire <= pkt_3_e_word_1337(31 downto 0);
    -- flow-through slice operator slice_1498_inst
    slice_1498_wire <= pkt_4_e_word_1342(31 downto 0);
    next_active_packet_1414_1350_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_active_packet_1414_1350_buf_req_0;
      next_active_packet_1414_1350_buf_ack_0<= wack(0);
      rreq(0) <= next_active_packet_1414_1350_buf_req_1;
      next_active_packet_1414_1350_buf_ack_1<= rack(0);
      next_active_packet_1414_1350_buf : InterlockBuffer generic map ( -- 
        name => "next_active_packet_1414_1350_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_active_packet_1414,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_active_packet_1414_1350_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_down_counter_1438_1326_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_down_counter_1438_1326_buf_req_0;
      next_down_counter_1438_1326_buf_ack_0<= wack(0);
      rreq(0) <= next_down_counter_1438_1326_buf_req_1;
      next_down_counter_1438_1326_buf_ack_1<= rack(0);
      next_down_counter_1438_1326_buf : InterlockBuffer generic map ( -- 
        name => "next_down_counter_1438_1326_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_down_counter_1438,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_down_counter_1438_1326_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_pkt_priority_1414_1354_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_pkt_priority_1414_1354_buf_req_0;
      next_pkt_priority_1414_1354_buf_ack_0<= wack(0);
      rreq(0) <= next_pkt_priority_1414_1354_buf_req_1;
      next_pkt_priority_1414_1354_buf_ack_1<= rack(0);
      next_pkt_priority_1414_1354_buf : InterlockBuffer generic map ( -- 
        name => "next_pkt_priority_1414_1354_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_pkt_priority_1414,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_pkt_priority_1414_1354_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1321_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1538_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1321_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1321_branch_req_0,
          ack0 => do_while_stmt_1321_branch_ack_0,
          ack1 => do_while_stmt_1321_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator AND_u1_u1_1426_inst
    process(OR_u1_u1_1422_wire, EQ_u8_u1_1425_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(OR_u1_u1_1422_wire, EQ_u8_u1_1425_wire, tmp_var);
      started_new_packet_1427 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_1359_inst
    process(pkt_1_e_word_1327) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_1_e_word_1327, konst_1358_wire_constant, tmp_var);
      p1_valid_1360 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_1364_inst
    process(pkt_2_e_word_1332) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_2_e_word_1332, konst_1363_wire_constant, tmp_var);
      p2_valid_1365 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_1369_inst
    process(pkt_3_e_word_1337) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_3_e_word_1337, konst_1368_wire_constant, tmp_var);
      p3_valid_1370 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u33_u1_1374_inst
    process(pkt_4_e_word_1342) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(pkt_4_e_word_1342, konst_1373_wire_constant, tmp_var);
      p4_valid_1375 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1379_inst
    process(active_packet_1347) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1347, konst_1378_wire_constant, tmp_var);
      EQ_u3_u1_1379_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1385_inst
    process(active_packet_1347) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1347, konst_1384_wire_constant, tmp_var);
      EQ_u3_u1_1385_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1392_inst
    process(active_packet_1347) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1347, konst_1391_wire_constant, tmp_var);
      EQ_u3_u1_1392_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1398_inst
    process(active_packet_1347) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(active_packet_1347, konst_1397_wire_constant, tmp_var);
      EQ_u3_u1_1398_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1444_inst
    process(next_active_packet_1414) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1414, konst_1443_wire_constant, tmp_var);
      EQ_u3_u1_1444_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1452_inst
    process(next_active_packet_1414) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1414, konst_1451_wire_constant, tmp_var);
      EQ_u3_u1_1452_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1460_inst
    process(next_active_packet_1414) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1414, konst_1459_wire_constant, tmp_var);
      EQ_u3_u1_1460_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1468_inst
    process(next_active_packet_1414) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1414, konst_1467_wire_constant, tmp_var);
      EQ_u3_u1_1468_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1474_inst
    process(next_active_packet_1414) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1414, konst_1473_wire_constant, tmp_var);
      EQ_u3_u1_1474_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1481_inst
    process(next_active_packet_1414) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1414, konst_1480_wire_constant, tmp_var);
      EQ_u3_u1_1481_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1489_inst
    process(next_active_packet_1414) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1414, konst_1488_wire_constant, tmp_var);
      EQ_u3_u1_1489_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1496_inst
    process(next_active_packet_1414) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1414, konst_1495_wire_constant, tmp_var);
      EQ_u3_u1_1496_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1507_inst
    process(next_active_packet_1414) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1414, konst_1506_wire_constant, tmp_var);
      EQ_u3_u1_1507_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1513_inst
    process(next_active_packet_1414) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1414, konst_1512_wire_constant, tmp_var);
      EQ_u3_u1_1513_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1520_inst
    process(next_active_packet_1414) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1414, konst_1519_wire_constant, tmp_var);
      EQ_u3_u1_1520_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1526_inst
    process(next_active_packet_1414) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_active_packet_1414, konst_1525_wire_constant, tmp_var);
      EQ_u3_u1_1526_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_1425_inst
    process(down_counter_1323) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(down_counter_1323, konst_1424_wire_constant, tmp_var);
      EQ_u8_u1_1425_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1441_inst
    process(p1_valid_1360) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_1360, tmp_var);
      NOT_u1_u1_1441_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1449_inst
    process(p2_valid_1365) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_1365, tmp_var);
      NOT_u1_u1_1449_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1457_inst
    process(p3_valid_1370) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_1370, tmp_var);
      NOT_u1_u1_1457_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1465_inst
    process(p4_valid_1375) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_1375, tmp_var);
      NOT_u1_u1_1465_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1389_inst
    process(MUX_1382_wire, MUX_1388_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1382_wire, MUX_1388_wire, tmp_var);
      OR_u1_u1_1389_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1402_inst
    process(MUX_1395_wire, MUX_1401_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1395_wire, MUX_1401_wire, tmp_var);
      OR_u1_u1_1402_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1403_inst
    process(OR_u1_u1_1389_wire, OR_u1_u1_1402_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1389_wire, OR_u1_u1_1402_wire, tmp_var);
      valid_active_pkt_word_read_1404 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1418_inst
    process(p1_valid_1360, p2_valid_1365) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(p1_valid_1360, p2_valid_1365, tmp_var);
      OR_u1_u1_1418_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1421_inst
    process(p3_valid_1370, p4_valid_1375) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(p3_valid_1370, p4_valid_1375, tmp_var);
      OR_u1_u1_1421_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1422_inst
    process(OR_u1_u1_1418_wire, OR_u1_u1_1421_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1418_wire, OR_u1_u1_1421_wire, tmp_var);
      OR_u1_u1_1422_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1445_inst
    process(NOT_u1_u1_1441_wire, EQ_u3_u1_1444_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1441_wire, EQ_u3_u1_1444_wire, tmp_var);
      read_from_1_1446 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1453_inst
    process(NOT_u1_u1_1449_wire, EQ_u3_u1_1452_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1449_wire, EQ_u3_u1_1452_wire, tmp_var);
      read_from_2_1454 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1461_inst
    process(NOT_u1_u1_1457_wire, EQ_u3_u1_1460_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1457_wire, EQ_u3_u1_1460_wire, tmp_var);
      read_from_3_1462 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1469_inst
    process(NOT_u1_u1_1465_wire, EQ_u3_u1_1468_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1465_wire, EQ_u3_u1_1468_wire, tmp_var);
      read_from_4_1470 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1517_inst
    process(MUX_1510_wire, MUX_1516_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1510_wire, MUX_1516_wire, tmp_var);
      OR_u1_u1_1517_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1530_inst
    process(MUX_1523_wire, MUX_1529_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1523_wire, MUX_1529_wire, tmp_var);
      OR_u1_u1_1530_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1531_inst
    process(OR_u1_u1_1517_wire, OR_u1_u1_1530_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1517_wire, OR_u1_u1_1530_wire, tmp_var);
      send_flag_1532 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1486_inst
    process(MUX_1478_wire, MUX_1485_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1478_wire, MUX_1485_wire, tmp_var);
      OR_u32_u32_1486_wire <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1501_inst
    process(MUX_1493_wire, MUX_1500_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1493_wire, MUX_1500_wire, tmp_var);
      OR_u32_u32_1501_wire <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1502_inst
    process(OR_u32_u32_1486_wire, OR_u32_u32_1501_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u32_u32_1486_wire, OR_u32_u32_1501_wire, tmp_var);
      data_to_out_1503 <= tmp_var; --
    end process;
    -- binary operator SUB_u8_u8_1434_inst
    process(down_counter_1323) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSub_proc(down_counter_1323, konst_1433_wire_constant, tmp_var);
      SUB_u8_u8_1434_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_noblock_obuf_1_4_1331_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_1_4_1331_inst_req_0;
      RPIPE_noblock_obuf_1_4_1331_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_1_4_1331_inst_req_1;
      RPIPE_noblock_obuf_1_4_1331_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_1_1446(0);
      RPIPE_noblock_obuf_1_4_1331_wire <= data_out(32 downto 0);
      noblock_obuf_1_4_read_0_gI: SplitGuardInterface generic map(name => "noblock_obuf_1_4_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_1_4_read_0: InputPortRevised -- 
        generic map ( name => "noblock_obuf_1_4_read_0", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_1_4_pipe_read_req(0),
          oack => noblock_obuf_1_4_pipe_read_ack(0),
          odata => noblock_obuf_1_4_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_noblock_obuf_2_4_1336_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_2_4_1336_inst_req_0;
      RPIPE_noblock_obuf_2_4_1336_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_2_4_1336_inst_req_1;
      RPIPE_noblock_obuf_2_4_1336_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_2_1454(0);
      RPIPE_noblock_obuf_2_4_1336_wire <= data_out(32 downto 0);
      noblock_obuf_2_4_read_1_gI: SplitGuardInterface generic map(name => "noblock_obuf_2_4_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_2_4_read_1: InputPortRevised -- 
        generic map ( name => "noblock_obuf_2_4_read_1", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_2_4_pipe_read_req(0),
          oack => noblock_obuf_2_4_pipe_read_ack(0),
          odata => noblock_obuf_2_4_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_noblock_obuf_3_4_1341_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_3_4_1341_inst_req_0;
      RPIPE_noblock_obuf_3_4_1341_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_3_4_1341_inst_req_1;
      RPIPE_noblock_obuf_3_4_1341_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_3_1462(0);
      RPIPE_noblock_obuf_3_4_1341_wire <= data_out(32 downto 0);
      noblock_obuf_3_4_read_2_gI: SplitGuardInterface generic map(name => "noblock_obuf_3_4_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_3_4_read_2: InputPortRevised -- 
        generic map ( name => "noblock_obuf_3_4_read_2", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_3_4_pipe_read_req(0),
          oack => noblock_obuf_3_4_pipe_read_ack(0),
          odata => noblock_obuf_3_4_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_noblock_obuf_4_4_1346_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_noblock_obuf_4_4_1346_inst_req_0;
      RPIPE_noblock_obuf_4_4_1346_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_noblock_obuf_4_4_1346_inst_req_1;
      RPIPE_noblock_obuf_4_4_1346_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_from_4_1470(0);
      RPIPE_noblock_obuf_4_4_1346_wire <= data_out(32 downto 0);
      noblock_obuf_4_4_read_3_gI: SplitGuardInterface generic map(name => "noblock_obuf_4_4_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      noblock_obuf_4_4_read_3: InputPortRevised -- 
        generic map ( name => "noblock_obuf_4_4_read_3", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => noblock_obuf_4_4_pipe_read_req(0),
          oack => noblock_obuf_4_4_pipe_read_ack(0),
          odata => noblock_obuf_4_4_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_out_data_4_1534_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_out_data_4_1534_inst_req_0;
      WPIPE_out_data_4_1534_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_out_data_4_1534_inst_req_1;
      WPIPE_out_data_4_1534_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_flag_1532(0);
      data_in <= data_to_out_1503;
      out_data_4_write_0_gI: SplitGuardInterface generic map(name => "out_data_4_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      out_data_4_write_0: OutputPortRevised -- 
        generic map ( name => "out_data_4", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => out_data_4_pipe_write_req(0),
          oack => out_data_4_pipe_write_ack(0),
          odata => out_data_4_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    volatile_operator_prioritySelect_3785: prioritySelect_Volatile port map(down_counter => down_counter_1323, active_packet => active_packet_1347, pkt_priority => pkt_priority_1351, p1_valid => p1_valid_1360, p2_valid => p2_valid_1365, p3_valid => p3_valid_1370, p4_valid => p4_valid_1375, next_active_packet => next_active_packet_1414, next_pkt_priority => next_pkt_priority_1414); 
    -- 
  end Block; -- data_path
  -- 
end outputPort_4_Daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity prioritySelect_Volatile is -- 
  port ( -- 
    down_counter : in  std_logic_vector(7 downto 0);
    active_packet : in  std_logic_vector(2 downto 0);
    pkt_priority : in  std_logic_vector(2 downto 0);
    p1_valid : in  std_logic_vector(0 downto 0);
    p2_valid : in  std_logic_vector(0 downto 0);
    p3_valid : in  std_logic_vector(0 downto 0);
    p4_valid : in  std_logic_vector(0 downto 0);
    next_active_packet : out  std_logic_vector(2 downto 0);
    next_pkt_priority : out  std_logic_vector(2 downto 0)-- 
  );
  -- 
end entity prioritySelect_Volatile;
architecture prioritySelect_Volatile_arch of prioritySelect_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(18-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal down_counter_buffer :  std_logic_vector(7 downto 0);
  signal active_packet_buffer :  std_logic_vector(2 downto 0);
  signal pkt_priority_buffer :  std_logic_vector(2 downto 0);
  signal p1_valid_buffer :  std_logic_vector(0 downto 0);
  signal p2_valid_buffer :  std_logic_vector(0 downto 0);
  signal p3_valid_buffer :  std_logic_vector(0 downto 0);
  signal p4_valid_buffer :  std_logic_vector(0 downto 0);
  -- output port buffer signals
  signal next_active_packet_buffer :  std_logic_vector(2 downto 0);
  signal next_pkt_priority_buffer :  std_logic_vector(2 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  down_counter_buffer <= down_counter;
  active_packet_buffer <= active_packet;
  pkt_priority_buffer <= pkt_priority;
  p1_valid_buffer <= p1_valid;
  p2_valid_buffer <= p2_valid;
  p3_valid_buffer <= p3_valid;
  p4_valid_buffer <= p4_valid;
  -- output handling  -------------------------------------------------------
  next_active_packet <= next_active_packet_buffer;
  next_pkt_priority <= next_pkt_priority_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_446_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_454_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_457_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_464_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_467_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_473_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_481_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_489_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_492_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_499_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_502_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_508_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_516_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_524_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_527_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_534_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_537_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_543_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_551_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_559_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_562_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_569_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_572_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_578_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_612_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_617_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_618_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_449_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_461_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_470_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_484_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_496_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_505_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_519_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_531_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_540_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_554_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_566_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_575_wire : std_logic_vector(0 downto 0);
    signal MUX_588_wire : std_logic_vector(2 downto 0);
    signal MUX_592_wire : std_logic_vector(2 downto 0);
    signal MUX_597_wire : std_logic_vector(2 downto 0);
    signal MUX_602_wire : std_logic_vector(2 downto 0);
    signal MUX_606_wire : std_logic_vector(2 downto 0);
    signal MUX_621_wire : std_logic_vector(2 downto 0);
    signal MUX_630_wire : std_logic_vector(2 downto 0);
    signal MUX_634_wire : std_logic_vector(2 downto 0);
    signal MUX_639_wire : std_logic_vector(2 downto 0);
    signal MUX_644_wire : std_logic_vector(2 downto 0);
    signal MUX_648_wire : std_logic_vector(2 downto 0);
    signal NOT_u1_u1_451_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_453_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_456_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_463_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_466_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_472_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_486_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_488_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_491_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_498_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_501_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_507_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_521_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_523_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_526_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_533_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_536_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_542_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_556_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_558_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_561_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_568_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_571_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_577_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_585_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_609_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_611_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_614_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_616_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_627_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_458_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_474_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_475_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_493_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_509_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_510_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_528_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_544_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_545_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_563_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_579_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_580_wire : std_logic_vector(0 downto 0);
    signal OR_u3_u3_593_wire : std_logic_vector(2 downto 0);
    signal OR_u3_u3_598_wire : std_logic_vector(2 downto 0);
    signal OR_u3_u3_607_wire : std_logic_vector(2 downto 0);
    signal OR_u3_u3_622_wire : std_logic_vector(2 downto 0);
    signal OR_u3_u3_635_wire : std_logic_vector(2 downto 0);
    signal OR_u3_u3_640_wire : std_logic_vector(2 downto 0);
    signal OR_u3_u3_649_wire : std_logic_vector(2 downto 0);
    signal d0_442 : std_logic_vector(0 downto 0);
    signal konst_440_wire_constant : std_logic_vector(7 downto 0);
    signal konst_448_wire_constant : std_logic_vector(2 downto 0);
    signal konst_460_wire_constant : std_logic_vector(2 downto 0);
    signal konst_469_wire_constant : std_logic_vector(2 downto 0);
    signal konst_483_wire_constant : std_logic_vector(2 downto 0);
    signal konst_495_wire_constant : std_logic_vector(2 downto 0);
    signal konst_504_wire_constant : std_logic_vector(2 downto 0);
    signal konst_518_wire_constant : std_logic_vector(2 downto 0);
    signal konst_530_wire_constant : std_logic_vector(2 downto 0);
    signal konst_539_wire_constant : std_logic_vector(2 downto 0);
    signal konst_553_wire_constant : std_logic_vector(2 downto 0);
    signal konst_565_wire_constant : std_logic_vector(2 downto 0);
    signal konst_574_wire_constant : std_logic_vector(2 downto 0);
    signal konst_587_wire_constant : std_logic_vector(2 downto 0);
    signal konst_590_wire_constant : std_logic_vector(2 downto 0);
    signal konst_591_wire_constant : std_logic_vector(2 downto 0);
    signal konst_595_wire_constant : std_logic_vector(2 downto 0);
    signal konst_596_wire_constant : std_logic_vector(2 downto 0);
    signal konst_600_wire_constant : std_logic_vector(2 downto 0);
    signal konst_601_wire_constant : std_logic_vector(2 downto 0);
    signal konst_604_wire_constant : std_logic_vector(2 downto 0);
    signal konst_605_wire_constant : std_logic_vector(2 downto 0);
    signal konst_620_wire_constant : std_logic_vector(2 downto 0);
    signal konst_629_wire_constant : std_logic_vector(2 downto 0);
    signal konst_632_wire_constant : std_logic_vector(2 downto 0);
    signal konst_633_wire_constant : std_logic_vector(2 downto 0);
    signal konst_637_wire_constant : std_logic_vector(2 downto 0);
    signal konst_638_wire_constant : std_logic_vector(2 downto 0);
    signal konst_642_wire_constant : std_logic_vector(2 downto 0);
    signal konst_643_wire_constant : std_logic_vector(2 downto 0);
    signal konst_646_wire_constant : std_logic_vector(2 downto 0);
    signal konst_647_wire_constant : std_logic_vector(2 downto 0);
    signal select_1_477 : std_logic_vector(0 downto 0);
    signal select_2_512 : std_logic_vector(0 downto 0);
    signal select_3_547 : std_logic_vector(0 downto 0);
    signal select_4_582 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    konst_440_wire_constant <= "00000000";
    konst_448_wire_constant <= "001";
    konst_460_wire_constant <= "011";
    konst_469_wire_constant <= "100";
    konst_483_wire_constant <= "010";
    konst_495_wire_constant <= "100";
    konst_504_wire_constant <= "001";
    konst_518_wire_constant <= "011";
    konst_530_wire_constant <= "001";
    konst_539_wire_constant <= "010";
    konst_553_wire_constant <= "100";
    konst_565_wire_constant <= "010";
    konst_574_wire_constant <= "011";
    konst_587_wire_constant <= "000";
    konst_590_wire_constant <= "001";
    konst_591_wire_constant <= "000";
    konst_595_wire_constant <= "010";
    konst_596_wire_constant <= "000";
    konst_600_wire_constant <= "011";
    konst_601_wire_constant <= "000";
    konst_604_wire_constant <= "100";
    konst_605_wire_constant <= "000";
    konst_620_wire_constant <= "000";
    konst_629_wire_constant <= "000";
    konst_632_wire_constant <= "010";
    konst_633_wire_constant <= "000";
    konst_637_wire_constant <= "011";
    konst_638_wire_constant <= "000";
    konst_642_wire_constant <= "100";
    konst_643_wire_constant <= "000";
    konst_646_wire_constant <= "001";
    konst_647_wire_constant <= "000";
    -- flow-through select operator MUX_588_inst
    MUX_588_wire <= active_packet_buffer when (NOT_u1_u1_585_wire(0) /=  '0') else konst_587_wire_constant;
    -- flow-through select operator MUX_592_inst
    MUX_592_wire <= konst_590_wire_constant when (select_1_477(0) /=  '0') else konst_591_wire_constant;
    -- flow-through select operator MUX_597_inst
    MUX_597_wire <= konst_595_wire_constant when (select_2_512(0) /=  '0') else konst_596_wire_constant;
    -- flow-through select operator MUX_602_inst
    MUX_602_wire <= konst_600_wire_constant when (select_3_547(0) /=  '0') else konst_601_wire_constant;
    -- flow-through select operator MUX_606_inst
    MUX_606_wire <= konst_604_wire_constant when (select_4_582(0) /=  '0') else konst_605_wire_constant;
    -- flow-through select operator MUX_621_inst
    MUX_621_wire <= active_packet_buffer when (AND_u1_u1_618_wire(0) /=  '0') else konst_620_wire_constant;
    -- flow-through select operator MUX_630_inst
    MUX_630_wire <= pkt_priority_buffer when (NOT_u1_u1_627_wire(0) /=  '0') else konst_629_wire_constant;
    -- flow-through select operator MUX_634_inst
    MUX_634_wire <= konst_632_wire_constant when (select_1_477(0) /=  '0') else konst_633_wire_constant;
    -- flow-through select operator MUX_639_inst
    MUX_639_wire <= konst_637_wire_constant when (select_2_512(0) /=  '0') else konst_638_wire_constant;
    -- flow-through select operator MUX_644_inst
    MUX_644_wire <= konst_642_wire_constant when (select_3_547(0) /=  '0') else konst_643_wire_constant;
    -- flow-through select operator MUX_648_inst
    MUX_648_wire <= konst_646_wire_constant when (select_4_582(0) /=  '0') else konst_647_wire_constant;
    -- binary operator AND_u1_u1_446_inst
    process(d0_442, p1_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(d0_442, p1_valid_buffer, tmp_var);
      AND_u1_u1_446_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_454_inst
    process(NOT_u1_u1_451_wire, NOT_u1_u1_453_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_451_wire, NOT_u1_u1_453_wire, tmp_var);
      AND_u1_u1_454_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_457_inst
    process(AND_u1_u1_454_wire, NOT_u1_u1_456_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_454_wire, NOT_u1_u1_456_wire, tmp_var);
      AND_u1_u1_457_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_464_inst
    process(EQ_u3_u1_461_wire, NOT_u1_u1_463_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u3_u1_461_wire, NOT_u1_u1_463_wire, tmp_var);
      AND_u1_u1_464_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_467_inst
    process(AND_u1_u1_464_wire, NOT_u1_u1_466_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_464_wire, NOT_u1_u1_466_wire, tmp_var);
      AND_u1_u1_467_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_473_inst
    process(EQ_u3_u1_470_wire, NOT_u1_u1_472_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u3_u1_470_wire, NOT_u1_u1_472_wire, tmp_var);
      AND_u1_u1_473_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_476_inst
    process(AND_u1_u1_446_wire, OR_u1_u1_475_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_446_wire, OR_u1_u1_475_wire, tmp_var);
      select_1_477 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_481_inst
    process(d0_442, p2_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(d0_442, p2_valid_buffer, tmp_var);
      AND_u1_u1_481_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_489_inst
    process(NOT_u1_u1_486_wire, NOT_u1_u1_488_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_486_wire, NOT_u1_u1_488_wire, tmp_var);
      AND_u1_u1_489_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_492_inst
    process(AND_u1_u1_489_wire, NOT_u1_u1_491_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_489_wire, NOT_u1_u1_491_wire, tmp_var);
      AND_u1_u1_492_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_499_inst
    process(EQ_u3_u1_496_wire, NOT_u1_u1_498_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u3_u1_496_wire, NOT_u1_u1_498_wire, tmp_var);
      AND_u1_u1_499_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_502_inst
    process(AND_u1_u1_499_wire, NOT_u1_u1_501_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_499_wire, NOT_u1_u1_501_wire, tmp_var);
      AND_u1_u1_502_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_508_inst
    process(EQ_u3_u1_505_wire, NOT_u1_u1_507_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u3_u1_505_wire, NOT_u1_u1_507_wire, tmp_var);
      AND_u1_u1_508_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_511_inst
    process(AND_u1_u1_481_wire, OR_u1_u1_510_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_481_wire, OR_u1_u1_510_wire, tmp_var);
      select_2_512 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_516_inst
    process(d0_442, p3_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(d0_442, p3_valid_buffer, tmp_var);
      AND_u1_u1_516_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_524_inst
    process(NOT_u1_u1_521_wire, NOT_u1_u1_523_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_521_wire, NOT_u1_u1_523_wire, tmp_var);
      AND_u1_u1_524_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_527_inst
    process(AND_u1_u1_524_wire, NOT_u1_u1_526_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_524_wire, NOT_u1_u1_526_wire, tmp_var);
      AND_u1_u1_527_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_534_inst
    process(EQ_u3_u1_531_wire, NOT_u1_u1_533_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u3_u1_531_wire, NOT_u1_u1_533_wire, tmp_var);
      AND_u1_u1_534_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_537_inst
    process(AND_u1_u1_534_wire, NOT_u1_u1_536_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_534_wire, NOT_u1_u1_536_wire, tmp_var);
      AND_u1_u1_537_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_543_inst
    process(EQ_u3_u1_540_wire, NOT_u1_u1_542_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u3_u1_540_wire, NOT_u1_u1_542_wire, tmp_var);
      AND_u1_u1_543_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_546_inst
    process(AND_u1_u1_516_wire, OR_u1_u1_545_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_516_wire, OR_u1_u1_545_wire, tmp_var);
      select_3_547 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_551_inst
    process(d0_442, p4_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(d0_442, p4_valid_buffer, tmp_var);
      AND_u1_u1_551_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_559_inst
    process(NOT_u1_u1_556_wire, NOT_u1_u1_558_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_556_wire, NOT_u1_u1_558_wire, tmp_var);
      AND_u1_u1_559_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_562_inst
    process(AND_u1_u1_559_wire, NOT_u1_u1_561_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_559_wire, NOT_u1_u1_561_wire, tmp_var);
      AND_u1_u1_562_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_569_inst
    process(EQ_u3_u1_566_wire, NOT_u1_u1_568_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u3_u1_566_wire, NOT_u1_u1_568_wire, tmp_var);
      AND_u1_u1_569_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_572_inst
    process(AND_u1_u1_569_wire, NOT_u1_u1_571_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_569_wire, NOT_u1_u1_571_wire, tmp_var);
      AND_u1_u1_572_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_578_inst
    process(EQ_u3_u1_575_wire, NOT_u1_u1_577_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u3_u1_575_wire, NOT_u1_u1_577_wire, tmp_var);
      AND_u1_u1_578_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_581_inst
    process(AND_u1_u1_551_wire, OR_u1_u1_580_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_551_wire, OR_u1_u1_580_wire, tmp_var);
      select_4_582 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_612_inst
    process(NOT_u1_u1_609_wire, NOT_u1_u1_611_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_609_wire, NOT_u1_u1_611_wire, tmp_var);
      AND_u1_u1_612_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_617_inst
    process(NOT_u1_u1_614_wire, NOT_u1_u1_616_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_614_wire, NOT_u1_u1_616_wire, tmp_var);
      AND_u1_u1_617_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_618_inst
    process(AND_u1_u1_612_wire, AND_u1_u1_617_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_612_wire, AND_u1_u1_617_wire, tmp_var);
      AND_u1_u1_618_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_449_inst
    process(pkt_priority_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(pkt_priority_buffer, konst_448_wire_constant, tmp_var);
      EQ_u3_u1_449_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_461_inst
    process(pkt_priority_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(pkt_priority_buffer, konst_460_wire_constant, tmp_var);
      EQ_u3_u1_461_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_470_inst
    process(pkt_priority_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(pkt_priority_buffer, konst_469_wire_constant, tmp_var);
      EQ_u3_u1_470_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_484_inst
    process(pkt_priority_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(pkt_priority_buffer, konst_483_wire_constant, tmp_var);
      EQ_u3_u1_484_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_496_inst
    process(pkt_priority_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(pkt_priority_buffer, konst_495_wire_constant, tmp_var);
      EQ_u3_u1_496_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_505_inst
    process(pkt_priority_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(pkt_priority_buffer, konst_504_wire_constant, tmp_var);
      EQ_u3_u1_505_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_519_inst
    process(pkt_priority_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(pkt_priority_buffer, konst_518_wire_constant, tmp_var);
      EQ_u3_u1_519_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_531_inst
    process(pkt_priority_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(pkt_priority_buffer, konst_530_wire_constant, tmp_var);
      EQ_u3_u1_531_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_540_inst
    process(pkt_priority_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(pkt_priority_buffer, konst_539_wire_constant, tmp_var);
      EQ_u3_u1_540_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_554_inst
    process(pkt_priority_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(pkt_priority_buffer, konst_553_wire_constant, tmp_var);
      EQ_u3_u1_554_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_566_inst
    process(pkt_priority_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(pkt_priority_buffer, konst_565_wire_constant, tmp_var);
      EQ_u3_u1_566_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_575_inst
    process(pkt_priority_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(pkt_priority_buffer, konst_574_wire_constant, tmp_var);
      EQ_u3_u1_575_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_441_inst
    process(down_counter_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(down_counter_buffer, konst_440_wire_constant, tmp_var);
      d0_442 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_451_inst
    process(p4_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_buffer, tmp_var);
      NOT_u1_u1_451_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_453_inst
    process(p2_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_buffer, tmp_var);
      NOT_u1_u1_453_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_456_inst
    process(p3_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_buffer, tmp_var);
      NOT_u1_u1_456_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_463_inst
    process(p3_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_buffer, tmp_var);
      NOT_u1_u1_463_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_466_inst
    process(p4_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_buffer, tmp_var);
      NOT_u1_u1_466_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_472_inst
    process(p4_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_buffer, tmp_var);
      NOT_u1_u1_472_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_486_inst
    process(p4_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_buffer, tmp_var);
      NOT_u1_u1_486_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_488_inst
    process(p1_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_buffer, tmp_var);
      NOT_u1_u1_488_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_491_inst
    process(p3_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_buffer, tmp_var);
      NOT_u1_u1_491_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_498_inst
    process(p4_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_buffer, tmp_var);
      NOT_u1_u1_498_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_501_inst
    process(p1_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_buffer, tmp_var);
      NOT_u1_u1_501_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_507_inst
    process(p1_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_buffer, tmp_var);
      NOT_u1_u1_507_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_521_inst
    process(p4_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p4_valid_buffer, tmp_var);
      NOT_u1_u1_521_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_523_inst
    process(p2_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_buffer, tmp_var);
      NOT_u1_u1_523_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_526_inst
    process(p1_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_buffer, tmp_var);
      NOT_u1_u1_526_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_533_inst
    process(p1_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_buffer, tmp_var);
      NOT_u1_u1_533_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_536_inst
    process(p2_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_buffer, tmp_var);
      NOT_u1_u1_536_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_542_inst
    process(p2_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_buffer, tmp_var);
      NOT_u1_u1_542_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_556_inst
    process(p1_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p1_valid_buffer, tmp_var);
      NOT_u1_u1_556_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_558_inst
    process(p2_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_buffer, tmp_var);
      NOT_u1_u1_558_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_561_inst
    process(p3_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_buffer, tmp_var);
      NOT_u1_u1_561_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_568_inst
    process(p2_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p2_valid_buffer, tmp_var);
      NOT_u1_u1_568_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_571_inst
    process(p3_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_buffer, tmp_var);
      NOT_u1_u1_571_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_577_inst
    process(p3_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", p3_valid_buffer, tmp_var);
      NOT_u1_u1_577_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_585_inst
    process(d0_442) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", d0_442, tmp_var);
      NOT_u1_u1_585_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_609_inst
    process(select_1_477) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", select_1_477, tmp_var);
      NOT_u1_u1_609_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_611_inst
    process(select_2_512) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", select_2_512, tmp_var);
      NOT_u1_u1_611_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_614_inst
    process(select_3_547) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", select_3_547, tmp_var);
      NOT_u1_u1_614_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_616_inst
    process(select_4_582) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", select_4_582, tmp_var);
      NOT_u1_u1_616_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_627_inst
    process(d0_442) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", d0_442, tmp_var);
      NOT_u1_u1_627_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_458_inst
    process(EQ_u3_u1_449_wire, AND_u1_u1_457_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u3_u1_449_wire, AND_u1_u1_457_wire, tmp_var);
      OR_u1_u1_458_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_474_inst
    process(AND_u1_u1_467_wire, AND_u1_u1_473_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_467_wire, AND_u1_u1_473_wire, tmp_var);
      OR_u1_u1_474_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_475_inst
    process(OR_u1_u1_458_wire, OR_u1_u1_474_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_458_wire, OR_u1_u1_474_wire, tmp_var);
      OR_u1_u1_475_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_493_inst
    process(EQ_u3_u1_484_wire, AND_u1_u1_492_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u3_u1_484_wire, AND_u1_u1_492_wire, tmp_var);
      OR_u1_u1_493_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_509_inst
    process(AND_u1_u1_502_wire, AND_u1_u1_508_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_502_wire, AND_u1_u1_508_wire, tmp_var);
      OR_u1_u1_509_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_510_inst
    process(OR_u1_u1_493_wire, OR_u1_u1_509_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_493_wire, OR_u1_u1_509_wire, tmp_var);
      OR_u1_u1_510_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_528_inst
    process(EQ_u3_u1_519_wire, AND_u1_u1_527_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u3_u1_519_wire, AND_u1_u1_527_wire, tmp_var);
      OR_u1_u1_528_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_544_inst
    process(AND_u1_u1_537_wire, AND_u1_u1_543_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_537_wire, AND_u1_u1_543_wire, tmp_var);
      OR_u1_u1_544_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_545_inst
    process(OR_u1_u1_528_wire, OR_u1_u1_544_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_528_wire, OR_u1_u1_544_wire, tmp_var);
      OR_u1_u1_545_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_563_inst
    process(EQ_u3_u1_554_wire, AND_u1_u1_562_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u3_u1_554_wire, AND_u1_u1_562_wire, tmp_var);
      OR_u1_u1_563_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_579_inst
    process(AND_u1_u1_572_wire, AND_u1_u1_578_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_572_wire, AND_u1_u1_578_wire, tmp_var);
      OR_u1_u1_579_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_580_inst
    process(OR_u1_u1_563_wire, OR_u1_u1_579_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_563_wire, OR_u1_u1_579_wire, tmp_var);
      OR_u1_u1_580_wire <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_593_inst
    process(MUX_588_wire, MUX_592_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_588_wire, MUX_592_wire, tmp_var);
      OR_u3_u3_593_wire <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_598_inst
    process(OR_u3_u3_593_wire, MUX_597_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u3_u3_593_wire, MUX_597_wire, tmp_var);
      OR_u3_u3_598_wire <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_607_inst
    process(MUX_602_wire, MUX_606_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_602_wire, MUX_606_wire, tmp_var);
      OR_u3_u3_607_wire <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_622_inst
    process(OR_u3_u3_607_wire, MUX_621_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u3_u3_607_wire, MUX_621_wire, tmp_var);
      OR_u3_u3_622_wire <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_623_inst
    process(OR_u3_u3_598_wire, OR_u3_u3_622_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u3_u3_598_wire, OR_u3_u3_622_wire, tmp_var);
      next_active_packet_buffer <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_635_inst
    process(MUX_630_wire, MUX_634_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_630_wire, MUX_634_wire, tmp_var);
      OR_u3_u3_635_wire <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_640_inst
    process(OR_u3_u3_635_wire, MUX_639_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u3_u3_635_wire, MUX_639_wire, tmp_var);
      OR_u3_u3_640_wire <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_649_inst
    process(MUX_644_wire, MUX_648_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_644_wire, MUX_648_wire, tmp_var);
      OR_u3_u3_649_wire <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_650_inst
    process(OR_u3_u3_640_wire, OR_u3_u3_649_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u3_u3_640_wire, OR_u3_u3_649_wire, tmp_var);
      next_pkt_priority_buffer <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end prioritySelect_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    in_data_1_pipe_write_data: in std_logic_vector(31 downto 0);
    in_data_1_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_1_pipe_write_ack : out std_logic_vector(0 downto 0);
    in_data_2_pipe_write_data: in std_logic_vector(31 downto 0);
    in_data_2_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_2_pipe_write_ack : out std_logic_vector(0 downto 0);
    in_data_3_pipe_write_data: in std_logic_vector(31 downto 0);
    in_data_3_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_3_pipe_write_ack : out std_logic_vector(0 downto 0);
    in_data_4_pipe_write_data: in std_logic_vector(31 downto 0);
    in_data_4_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_4_pipe_write_ack : out std_logic_vector(0 downto 0);
    out_data_1_pipe_read_data: out std_logic_vector(31 downto 0);
    out_data_1_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_1_pipe_read_ack : out std_logic_vector(0 downto 0);
    out_data_2_pipe_read_data: out std_logic_vector(31 downto 0);
    out_data_2_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_2_pipe_read_ack : out std_logic_vector(0 downto 0);
    out_data_3_pipe_read_data: out std_logic_vector(31 downto 0);
    out_data_3_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_3_pipe_read_ack : out std_logic_vector(0 downto 0);
    out_data_4_pipe_read_data: out std_logic_vector(31 downto 0);
    out_data_4_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_4_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- declarations related to module inputPort_1_Daemon
  component inputPort_1_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      in_data_1_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_1_pipe_read_data : in   std_logic_vector(31 downto 0);
      noblock_obuf_1_3_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_3_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_1_4_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_4_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_1_1_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_1_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_1_2_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_2_pipe_write_data : out  std_logic_vector(32 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module inputPort_1_Daemon
  signal inputPort_1_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal inputPort_1_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal inputPort_1_Daemon_start_req : std_logic;
  signal inputPort_1_Daemon_start_ack : std_logic;
  signal inputPort_1_Daemon_fin_req   : std_logic;
  signal inputPort_1_Daemon_fin_ack : std_logic;
  -- declarations related to module inputPort_2_Daemon
  component inputPort_2_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      in_data_2_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_2_pipe_read_data : in   std_logic_vector(31 downto 0);
      noblock_obuf_2_1_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_1_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_2_2_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_2_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_2_3_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_3_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_2_4_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_4_pipe_write_data : out  std_logic_vector(32 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module inputPort_2_Daemon
  signal inputPort_2_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal inputPort_2_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal inputPort_2_Daemon_start_req : std_logic;
  signal inputPort_2_Daemon_start_ack : std_logic;
  signal inputPort_2_Daemon_fin_req   : std_logic;
  signal inputPort_2_Daemon_fin_ack : std_logic;
  -- declarations related to module inputPort_3_Daemon
  component inputPort_3_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      in_data_3_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_3_pipe_read_data : in   std_logic_vector(31 downto 0);
      noblock_obuf_3_2_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_2_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_3_3_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_3_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_3_4_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_4_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_3_1_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_1_pipe_write_data : out  std_logic_vector(32 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module inputPort_3_Daemon
  signal inputPort_3_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal inputPort_3_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal inputPort_3_Daemon_start_req : std_logic;
  signal inputPort_3_Daemon_start_ack : std_logic;
  signal inputPort_3_Daemon_fin_req   : std_logic;
  signal inputPort_3_Daemon_fin_ack : std_logic;
  -- declarations related to module inputPort_4_Daemon
  component inputPort_4_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      in_data_4_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_4_pipe_read_data : in   std_logic_vector(31 downto 0);
      noblock_obuf_4_1_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_1_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_4_2_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_2_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_4_3_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_3_pipe_write_data : out  std_logic_vector(32 downto 0);
      noblock_obuf_4_4_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_4_pipe_write_data : out  std_logic_vector(32 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module inputPort_4_Daemon
  signal inputPort_4_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal inputPort_4_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal inputPort_4_Daemon_start_req : std_logic;
  signal inputPort_4_Daemon_start_ack : std_logic;
  signal inputPort_4_Daemon_fin_req   : std_logic;
  signal inputPort_4_Daemon_fin_ack : std_logic;
  -- declarations related to module outputPort_1_Daemon
  component outputPort_1_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      noblock_obuf_4_1_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_1_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_2_1_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_1_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_1_1_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_1_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_3_1_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_1_pipe_read_data : in   std_logic_vector(32 downto 0);
      out_data_1_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_1_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module outputPort_1_Daemon
  signal outputPort_1_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal outputPort_1_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal outputPort_1_Daemon_start_req : std_logic;
  signal outputPort_1_Daemon_start_ack : std_logic;
  signal outputPort_1_Daemon_fin_req   : std_logic;
  signal outputPort_1_Daemon_fin_ack : std_logic;
  -- declarations related to module outputPort_2_Daemon
  component outputPort_2_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      noblock_obuf_1_2_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_2_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_3_2_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_2_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_4_2_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_2_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_2_2_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_2_pipe_read_data : in   std_logic_vector(32 downto 0);
      out_data_2_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_2_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module outputPort_2_Daemon
  signal outputPort_2_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal outputPort_2_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal outputPort_2_Daemon_start_req : std_logic;
  signal outputPort_2_Daemon_start_ack : std_logic;
  signal outputPort_2_Daemon_fin_req   : std_logic;
  signal outputPort_2_Daemon_fin_ack : std_logic;
  -- declarations related to module outputPort_3_Daemon
  component outputPort_3_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      noblock_obuf_1_3_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_3_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_3_3_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_3_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_4_3_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_3_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_2_3_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_3_pipe_read_data : in   std_logic_vector(32 downto 0);
      out_data_3_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_3_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module outputPort_3_Daemon
  signal outputPort_3_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal outputPort_3_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal outputPort_3_Daemon_start_req : std_logic;
  signal outputPort_3_Daemon_start_ack : std_logic;
  signal outputPort_3_Daemon_fin_req   : std_logic;
  signal outputPort_3_Daemon_fin_ack : std_logic;
  -- declarations related to module outputPort_4_Daemon
  component outputPort_4_Daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      noblock_obuf_1_4_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_1_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_1_4_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_3_4_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_3_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_3_4_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_2_4_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_2_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_2_4_pipe_read_data : in   std_logic_vector(32 downto 0);
      noblock_obuf_4_4_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_obuf_4_4_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_obuf_4_4_pipe_read_data : in   std_logic_vector(32 downto 0);
      out_data_4_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_4_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module outputPort_4_Daemon
  signal outputPort_4_Daemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal outputPort_4_Daemon_tag_out   : std_logic_vector(1 downto 0);
  signal outputPort_4_Daemon_start_req : std_logic;
  signal outputPort_4_Daemon_start_ack : std_logic;
  signal outputPort_4_Daemon_fin_req   : std_logic;
  signal outputPort_4_Daemon_fin_ack : std_logic;
  -- declarations related to module prioritySelect
  -- aggregate signals for read from pipe in_data_1
  signal in_data_1_pipe_read_data: std_logic_vector(31 downto 0);
  signal in_data_1_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_data_2
  signal in_data_2_pipe_read_data: std_logic_vector(31 downto 0);
  signal in_data_2_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_data_3
  signal in_data_3_pipe_read_data: std_logic_vector(31 downto 0);
  signal in_data_3_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_data_4
  signal in_data_4_pipe_read_data: std_logic_vector(31 downto 0);
  signal in_data_4_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_4_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_1_1
  signal noblock_obuf_1_1_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_1_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_1_1
  signal noblock_obuf_1_1_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_1_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_1_2
  signal noblock_obuf_1_2_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_2_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_1_2
  signal noblock_obuf_1_2_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_2_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_1_3
  signal noblock_obuf_1_3_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_3_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_1_3
  signal noblock_obuf_1_3_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_3_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_1_4
  signal noblock_obuf_1_4_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_4_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_4_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_1_4
  signal noblock_obuf_1_4_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_1_4_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_1_4_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_2_1
  signal noblock_obuf_2_1_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_1_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_2_1
  signal noblock_obuf_2_1_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_1_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_2_2
  signal noblock_obuf_2_2_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_2_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_2_2
  signal noblock_obuf_2_2_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_2_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_2_3
  signal noblock_obuf_2_3_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_3_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_2_3
  signal noblock_obuf_2_3_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_3_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_2_4
  signal noblock_obuf_2_4_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_4_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_4_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_2_4
  signal noblock_obuf_2_4_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_2_4_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_2_4_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_3_1
  signal noblock_obuf_3_1_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_1_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_3_1
  signal noblock_obuf_3_1_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_1_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_3_2
  signal noblock_obuf_3_2_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_2_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_3_2
  signal noblock_obuf_3_2_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_2_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_3_3
  signal noblock_obuf_3_3_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_3_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_3_3
  signal noblock_obuf_3_3_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_3_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_3_4
  signal noblock_obuf_3_4_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_4_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_4_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_3_4
  signal noblock_obuf_3_4_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_3_4_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_3_4_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_4_1
  signal noblock_obuf_4_1_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_1_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_4_1
  signal noblock_obuf_4_1_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_1_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_4_2
  signal noblock_obuf_4_2_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_2_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_4_2
  signal noblock_obuf_4_2_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_2_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_4_3
  signal noblock_obuf_4_3_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_3_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_4_3
  signal noblock_obuf_4_3_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_3_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe noblock_obuf_4_4
  signal noblock_obuf_4_4_pipe_write_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_4_pipe_write_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_4_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe noblock_obuf_4_4
  signal noblock_obuf_4_4_pipe_read_data: std_logic_vector(32 downto 0);
  signal noblock_obuf_4_4_pipe_read_req: std_logic_vector(0 downto 0);
  signal noblock_obuf_4_4_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data_1
  signal out_data_1_pipe_write_data: std_logic_vector(31 downto 0);
  signal out_data_1_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data_2
  signal out_data_2_pipe_write_data: std_logic_vector(31 downto 0);
  signal out_data_2_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data_3
  signal out_data_3_pipe_write_data: std_logic_vector(31 downto 0);
  signal out_data_3_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data_4
  signal out_data_4_pipe_write_data: std_logic_vector(31 downto 0);
  signal out_data_4_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_4_pipe_write_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module inputPort_1_Daemon
  inputPort_1_Daemon_instance:inputPort_1_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => inputPort_1_Daemon_start_req,
      start_ack => inputPort_1_Daemon_start_ack,
      fin_req => inputPort_1_Daemon_fin_req,
      fin_ack => inputPort_1_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      in_data_1_pipe_read_req => in_data_1_pipe_read_req(0 downto 0),
      in_data_1_pipe_read_ack => in_data_1_pipe_read_ack(0 downto 0),
      in_data_1_pipe_read_data => in_data_1_pipe_read_data(31 downto 0),
      noblock_obuf_1_3_pipe_write_req => noblock_obuf_1_3_pipe_write_req(0 downto 0),
      noblock_obuf_1_3_pipe_write_ack => noblock_obuf_1_3_pipe_write_ack(0 downto 0),
      noblock_obuf_1_3_pipe_write_data => noblock_obuf_1_3_pipe_write_data(32 downto 0),
      noblock_obuf_1_4_pipe_write_req => noblock_obuf_1_4_pipe_write_req(0 downto 0),
      noblock_obuf_1_4_pipe_write_ack => noblock_obuf_1_4_pipe_write_ack(0 downto 0),
      noblock_obuf_1_4_pipe_write_data => noblock_obuf_1_4_pipe_write_data(32 downto 0),
      noblock_obuf_1_1_pipe_write_req => noblock_obuf_1_1_pipe_write_req(0 downto 0),
      noblock_obuf_1_1_pipe_write_ack => noblock_obuf_1_1_pipe_write_ack(0 downto 0),
      noblock_obuf_1_1_pipe_write_data => noblock_obuf_1_1_pipe_write_data(32 downto 0),
      noblock_obuf_1_2_pipe_write_req => noblock_obuf_1_2_pipe_write_req(0 downto 0),
      noblock_obuf_1_2_pipe_write_ack => noblock_obuf_1_2_pipe_write_ack(0 downto 0),
      noblock_obuf_1_2_pipe_write_data => noblock_obuf_1_2_pipe_write_data(32 downto 0),
      tag_in => inputPort_1_Daemon_tag_in,
      tag_out => inputPort_1_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  inputPort_1_Daemon_tag_in <= (others => '0');
  inputPort_1_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => inputPort_1_Daemon_start_req, start_ack => inputPort_1_Daemon_start_ack,  fin_req => inputPort_1_Daemon_fin_req,  fin_ack => inputPort_1_Daemon_fin_ack);
  -- module inputPort_2_Daemon
  inputPort_2_Daemon_instance:inputPort_2_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => inputPort_2_Daemon_start_req,
      start_ack => inputPort_2_Daemon_start_ack,
      fin_req => inputPort_2_Daemon_fin_req,
      fin_ack => inputPort_2_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      in_data_2_pipe_read_req => in_data_2_pipe_read_req(0 downto 0),
      in_data_2_pipe_read_ack => in_data_2_pipe_read_ack(0 downto 0),
      in_data_2_pipe_read_data => in_data_2_pipe_read_data(31 downto 0),
      noblock_obuf_2_1_pipe_write_req => noblock_obuf_2_1_pipe_write_req(0 downto 0),
      noblock_obuf_2_1_pipe_write_ack => noblock_obuf_2_1_pipe_write_ack(0 downto 0),
      noblock_obuf_2_1_pipe_write_data => noblock_obuf_2_1_pipe_write_data(32 downto 0),
      noblock_obuf_2_2_pipe_write_req => noblock_obuf_2_2_pipe_write_req(0 downto 0),
      noblock_obuf_2_2_pipe_write_ack => noblock_obuf_2_2_pipe_write_ack(0 downto 0),
      noblock_obuf_2_2_pipe_write_data => noblock_obuf_2_2_pipe_write_data(32 downto 0),
      noblock_obuf_2_3_pipe_write_req => noblock_obuf_2_3_pipe_write_req(0 downto 0),
      noblock_obuf_2_3_pipe_write_ack => noblock_obuf_2_3_pipe_write_ack(0 downto 0),
      noblock_obuf_2_3_pipe_write_data => noblock_obuf_2_3_pipe_write_data(32 downto 0),
      noblock_obuf_2_4_pipe_write_req => noblock_obuf_2_4_pipe_write_req(0 downto 0),
      noblock_obuf_2_4_pipe_write_ack => noblock_obuf_2_4_pipe_write_ack(0 downto 0),
      noblock_obuf_2_4_pipe_write_data => noblock_obuf_2_4_pipe_write_data(32 downto 0),
      tag_in => inputPort_2_Daemon_tag_in,
      tag_out => inputPort_2_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  inputPort_2_Daemon_tag_in <= (others => '0');
  inputPort_2_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => inputPort_2_Daemon_start_req, start_ack => inputPort_2_Daemon_start_ack,  fin_req => inputPort_2_Daemon_fin_req,  fin_ack => inputPort_2_Daemon_fin_ack);
  -- module inputPort_3_Daemon
  inputPort_3_Daemon_instance:inputPort_3_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => inputPort_3_Daemon_start_req,
      start_ack => inputPort_3_Daemon_start_ack,
      fin_req => inputPort_3_Daemon_fin_req,
      fin_ack => inputPort_3_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      in_data_3_pipe_read_req => in_data_3_pipe_read_req(0 downto 0),
      in_data_3_pipe_read_ack => in_data_3_pipe_read_ack(0 downto 0),
      in_data_3_pipe_read_data => in_data_3_pipe_read_data(31 downto 0),
      noblock_obuf_3_2_pipe_write_req => noblock_obuf_3_2_pipe_write_req(0 downto 0),
      noblock_obuf_3_2_pipe_write_ack => noblock_obuf_3_2_pipe_write_ack(0 downto 0),
      noblock_obuf_3_2_pipe_write_data => noblock_obuf_3_2_pipe_write_data(32 downto 0),
      noblock_obuf_3_3_pipe_write_req => noblock_obuf_3_3_pipe_write_req(0 downto 0),
      noblock_obuf_3_3_pipe_write_ack => noblock_obuf_3_3_pipe_write_ack(0 downto 0),
      noblock_obuf_3_3_pipe_write_data => noblock_obuf_3_3_pipe_write_data(32 downto 0),
      noblock_obuf_3_4_pipe_write_req => noblock_obuf_3_4_pipe_write_req(0 downto 0),
      noblock_obuf_3_4_pipe_write_ack => noblock_obuf_3_4_pipe_write_ack(0 downto 0),
      noblock_obuf_3_4_pipe_write_data => noblock_obuf_3_4_pipe_write_data(32 downto 0),
      noblock_obuf_3_1_pipe_write_req => noblock_obuf_3_1_pipe_write_req(0 downto 0),
      noblock_obuf_3_1_pipe_write_ack => noblock_obuf_3_1_pipe_write_ack(0 downto 0),
      noblock_obuf_3_1_pipe_write_data => noblock_obuf_3_1_pipe_write_data(32 downto 0),
      tag_in => inputPort_3_Daemon_tag_in,
      tag_out => inputPort_3_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  inputPort_3_Daemon_tag_in <= (others => '0');
  inputPort_3_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => inputPort_3_Daemon_start_req, start_ack => inputPort_3_Daemon_start_ack,  fin_req => inputPort_3_Daemon_fin_req,  fin_ack => inputPort_3_Daemon_fin_ack);
  -- module inputPort_4_Daemon
  inputPort_4_Daemon_instance:inputPort_4_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => inputPort_4_Daemon_start_req,
      start_ack => inputPort_4_Daemon_start_ack,
      fin_req => inputPort_4_Daemon_fin_req,
      fin_ack => inputPort_4_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      in_data_4_pipe_read_req => in_data_4_pipe_read_req(0 downto 0),
      in_data_4_pipe_read_ack => in_data_4_pipe_read_ack(0 downto 0),
      in_data_4_pipe_read_data => in_data_4_pipe_read_data(31 downto 0),
      noblock_obuf_4_1_pipe_write_req => noblock_obuf_4_1_pipe_write_req(0 downto 0),
      noblock_obuf_4_1_pipe_write_ack => noblock_obuf_4_1_pipe_write_ack(0 downto 0),
      noblock_obuf_4_1_pipe_write_data => noblock_obuf_4_1_pipe_write_data(32 downto 0),
      noblock_obuf_4_2_pipe_write_req => noblock_obuf_4_2_pipe_write_req(0 downto 0),
      noblock_obuf_4_2_pipe_write_ack => noblock_obuf_4_2_pipe_write_ack(0 downto 0),
      noblock_obuf_4_2_pipe_write_data => noblock_obuf_4_2_pipe_write_data(32 downto 0),
      noblock_obuf_4_3_pipe_write_req => noblock_obuf_4_3_pipe_write_req(0 downto 0),
      noblock_obuf_4_3_pipe_write_ack => noblock_obuf_4_3_pipe_write_ack(0 downto 0),
      noblock_obuf_4_3_pipe_write_data => noblock_obuf_4_3_pipe_write_data(32 downto 0),
      noblock_obuf_4_4_pipe_write_req => noblock_obuf_4_4_pipe_write_req(0 downto 0),
      noblock_obuf_4_4_pipe_write_ack => noblock_obuf_4_4_pipe_write_ack(0 downto 0),
      noblock_obuf_4_4_pipe_write_data => noblock_obuf_4_4_pipe_write_data(32 downto 0),
      tag_in => inputPort_4_Daemon_tag_in,
      tag_out => inputPort_4_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  inputPort_4_Daemon_tag_in <= (others => '0');
  inputPort_4_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => inputPort_4_Daemon_start_req, start_ack => inputPort_4_Daemon_start_ack,  fin_req => inputPort_4_Daemon_fin_req,  fin_ack => inputPort_4_Daemon_fin_ack);
  -- module outputPort_1_Daemon
  outputPort_1_Daemon_instance:outputPort_1_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => outputPort_1_Daemon_start_req,
      start_ack => outputPort_1_Daemon_start_ack,
      fin_req => outputPort_1_Daemon_fin_req,
      fin_ack => outputPort_1_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      noblock_obuf_4_1_pipe_read_req => noblock_obuf_4_1_pipe_read_req(0 downto 0),
      noblock_obuf_4_1_pipe_read_ack => noblock_obuf_4_1_pipe_read_ack(0 downto 0),
      noblock_obuf_4_1_pipe_read_data => noblock_obuf_4_1_pipe_read_data(32 downto 0),
      noblock_obuf_2_1_pipe_read_req => noblock_obuf_2_1_pipe_read_req(0 downto 0),
      noblock_obuf_2_1_pipe_read_ack => noblock_obuf_2_1_pipe_read_ack(0 downto 0),
      noblock_obuf_2_1_pipe_read_data => noblock_obuf_2_1_pipe_read_data(32 downto 0),
      noblock_obuf_1_1_pipe_read_req => noblock_obuf_1_1_pipe_read_req(0 downto 0),
      noblock_obuf_1_1_pipe_read_ack => noblock_obuf_1_1_pipe_read_ack(0 downto 0),
      noblock_obuf_1_1_pipe_read_data => noblock_obuf_1_1_pipe_read_data(32 downto 0),
      noblock_obuf_3_1_pipe_read_req => noblock_obuf_3_1_pipe_read_req(0 downto 0),
      noblock_obuf_3_1_pipe_read_ack => noblock_obuf_3_1_pipe_read_ack(0 downto 0),
      noblock_obuf_3_1_pipe_read_data => noblock_obuf_3_1_pipe_read_data(32 downto 0),
      out_data_1_pipe_write_req => out_data_1_pipe_write_req(0 downto 0),
      out_data_1_pipe_write_ack => out_data_1_pipe_write_ack(0 downto 0),
      out_data_1_pipe_write_data => out_data_1_pipe_write_data(31 downto 0),
      tag_in => outputPort_1_Daemon_tag_in,
      tag_out => outputPort_1_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  outputPort_1_Daemon_tag_in <= (others => '0');
  outputPort_1_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => outputPort_1_Daemon_start_req, start_ack => outputPort_1_Daemon_start_ack,  fin_req => outputPort_1_Daemon_fin_req,  fin_ack => outputPort_1_Daemon_fin_ack);
  -- module outputPort_2_Daemon
  outputPort_2_Daemon_instance:outputPort_2_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => outputPort_2_Daemon_start_req,
      start_ack => outputPort_2_Daemon_start_ack,
      fin_req => outputPort_2_Daemon_fin_req,
      fin_ack => outputPort_2_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      noblock_obuf_1_2_pipe_read_req => noblock_obuf_1_2_pipe_read_req(0 downto 0),
      noblock_obuf_1_2_pipe_read_ack => noblock_obuf_1_2_pipe_read_ack(0 downto 0),
      noblock_obuf_1_2_pipe_read_data => noblock_obuf_1_2_pipe_read_data(32 downto 0),
      noblock_obuf_3_2_pipe_read_req => noblock_obuf_3_2_pipe_read_req(0 downto 0),
      noblock_obuf_3_2_pipe_read_ack => noblock_obuf_3_2_pipe_read_ack(0 downto 0),
      noblock_obuf_3_2_pipe_read_data => noblock_obuf_3_2_pipe_read_data(32 downto 0),
      noblock_obuf_4_2_pipe_read_req => noblock_obuf_4_2_pipe_read_req(0 downto 0),
      noblock_obuf_4_2_pipe_read_ack => noblock_obuf_4_2_pipe_read_ack(0 downto 0),
      noblock_obuf_4_2_pipe_read_data => noblock_obuf_4_2_pipe_read_data(32 downto 0),
      noblock_obuf_2_2_pipe_read_req => noblock_obuf_2_2_pipe_read_req(0 downto 0),
      noblock_obuf_2_2_pipe_read_ack => noblock_obuf_2_2_pipe_read_ack(0 downto 0),
      noblock_obuf_2_2_pipe_read_data => noblock_obuf_2_2_pipe_read_data(32 downto 0),
      out_data_2_pipe_write_req => out_data_2_pipe_write_req(0 downto 0),
      out_data_2_pipe_write_ack => out_data_2_pipe_write_ack(0 downto 0),
      out_data_2_pipe_write_data => out_data_2_pipe_write_data(31 downto 0),
      tag_in => outputPort_2_Daemon_tag_in,
      tag_out => outputPort_2_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  outputPort_2_Daemon_tag_in <= (others => '0');
  outputPort_2_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => outputPort_2_Daemon_start_req, start_ack => outputPort_2_Daemon_start_ack,  fin_req => outputPort_2_Daemon_fin_req,  fin_ack => outputPort_2_Daemon_fin_ack);
  -- module outputPort_3_Daemon
  outputPort_3_Daemon_instance:outputPort_3_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => outputPort_3_Daemon_start_req,
      start_ack => outputPort_3_Daemon_start_ack,
      fin_req => outputPort_3_Daemon_fin_req,
      fin_ack => outputPort_3_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      noblock_obuf_1_3_pipe_read_req => noblock_obuf_1_3_pipe_read_req(0 downto 0),
      noblock_obuf_1_3_pipe_read_ack => noblock_obuf_1_3_pipe_read_ack(0 downto 0),
      noblock_obuf_1_3_pipe_read_data => noblock_obuf_1_3_pipe_read_data(32 downto 0),
      noblock_obuf_3_3_pipe_read_req => noblock_obuf_3_3_pipe_read_req(0 downto 0),
      noblock_obuf_3_3_pipe_read_ack => noblock_obuf_3_3_pipe_read_ack(0 downto 0),
      noblock_obuf_3_3_pipe_read_data => noblock_obuf_3_3_pipe_read_data(32 downto 0),
      noblock_obuf_4_3_pipe_read_req => noblock_obuf_4_3_pipe_read_req(0 downto 0),
      noblock_obuf_4_3_pipe_read_ack => noblock_obuf_4_3_pipe_read_ack(0 downto 0),
      noblock_obuf_4_3_pipe_read_data => noblock_obuf_4_3_pipe_read_data(32 downto 0),
      noblock_obuf_2_3_pipe_read_req => noblock_obuf_2_3_pipe_read_req(0 downto 0),
      noblock_obuf_2_3_pipe_read_ack => noblock_obuf_2_3_pipe_read_ack(0 downto 0),
      noblock_obuf_2_3_pipe_read_data => noblock_obuf_2_3_pipe_read_data(32 downto 0),
      out_data_3_pipe_write_req => out_data_3_pipe_write_req(0 downto 0),
      out_data_3_pipe_write_ack => out_data_3_pipe_write_ack(0 downto 0),
      out_data_3_pipe_write_data => out_data_3_pipe_write_data(31 downto 0),
      tag_in => outputPort_3_Daemon_tag_in,
      tag_out => outputPort_3_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  outputPort_3_Daemon_tag_in <= (others => '0');
  outputPort_3_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => outputPort_3_Daemon_start_req, start_ack => outputPort_3_Daemon_start_ack,  fin_req => outputPort_3_Daemon_fin_req,  fin_ack => outputPort_3_Daemon_fin_ack);
  -- module outputPort_4_Daemon
  outputPort_4_Daemon_instance:outputPort_4_Daemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => outputPort_4_Daemon_start_req,
      start_ack => outputPort_4_Daemon_start_ack,
      fin_req => outputPort_4_Daemon_fin_req,
      fin_ack => outputPort_4_Daemon_fin_ack,
      clk => clk,
      reset => reset,
      noblock_obuf_1_4_pipe_read_req => noblock_obuf_1_4_pipe_read_req(0 downto 0),
      noblock_obuf_1_4_pipe_read_ack => noblock_obuf_1_4_pipe_read_ack(0 downto 0),
      noblock_obuf_1_4_pipe_read_data => noblock_obuf_1_4_pipe_read_data(32 downto 0),
      noblock_obuf_3_4_pipe_read_req => noblock_obuf_3_4_pipe_read_req(0 downto 0),
      noblock_obuf_3_4_pipe_read_ack => noblock_obuf_3_4_pipe_read_ack(0 downto 0),
      noblock_obuf_3_4_pipe_read_data => noblock_obuf_3_4_pipe_read_data(32 downto 0),
      noblock_obuf_2_4_pipe_read_req => noblock_obuf_2_4_pipe_read_req(0 downto 0),
      noblock_obuf_2_4_pipe_read_ack => noblock_obuf_2_4_pipe_read_ack(0 downto 0),
      noblock_obuf_2_4_pipe_read_data => noblock_obuf_2_4_pipe_read_data(32 downto 0),
      noblock_obuf_4_4_pipe_read_req => noblock_obuf_4_4_pipe_read_req(0 downto 0),
      noblock_obuf_4_4_pipe_read_ack => noblock_obuf_4_4_pipe_read_ack(0 downto 0),
      noblock_obuf_4_4_pipe_read_data => noblock_obuf_4_4_pipe_read_data(32 downto 0),
      out_data_4_pipe_write_req => out_data_4_pipe_write_req(0 downto 0),
      out_data_4_pipe_write_ack => out_data_4_pipe_write_ack(0 downto 0),
      out_data_4_pipe_write_data => out_data_4_pipe_write_data(31 downto 0),
      tag_in => outputPort_4_Daemon_tag_in,
      tag_out => outputPort_4_Daemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  outputPort_4_Daemon_tag_in <= (others => '0');
  outputPort_4_Daemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => outputPort_4_Daemon_start_req, start_ack => outputPort_4_Daemon_start_ack,  fin_req => outputPort_4_Daemon_fin_req,  fin_ack => outputPort_4_Daemon_fin_ack);
  in_data_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe in_data_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => in_data_1_pipe_read_req,
      read_ack => in_data_1_pipe_read_ack,
      read_data => in_data_1_pipe_read_data,
      write_req => in_data_1_pipe_write_req,
      write_ack => in_data_1_pipe_write_ack,
      write_data => in_data_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  in_data_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe in_data_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => in_data_2_pipe_read_req,
      read_ack => in_data_2_pipe_read_ack,
      read_data => in_data_2_pipe_read_data,
      write_req => in_data_2_pipe_write_req,
      write_ack => in_data_2_pipe_write_ack,
      write_data => in_data_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  in_data_3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe in_data_3",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => in_data_3_pipe_read_req,
      read_ack => in_data_3_pipe_read_ack,
      read_data => in_data_3_pipe_read_data,
      write_req => in_data_3_pipe_write_req,
      write_ack => in_data_3_pipe_write_ack,
      write_data => in_data_3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  in_data_4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe in_data_4",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => in_data_4_pipe_read_req,
      read_ack => in_data_4_pipe_read_ack,
      read_data => in_data_4_pipe_read_data,
      write_req => in_data_4_pipe_write_req,
      write_ack => in_data_4_pipe_write_ack,
      write_data => in_data_4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_1_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_1_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_1_1_pipe_read_req,
      read_ack => noblock_obuf_1_1_pipe_read_ack,
      read_data => noblock_obuf_1_1_pipe_read_data,
      write_req => noblock_obuf_1_1_pipe_write_req,
      write_ack => noblock_obuf_1_1_pipe_write_ack,
      write_data => noblock_obuf_1_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_1_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_1_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_1_2_pipe_read_req,
      read_ack => noblock_obuf_1_2_pipe_read_ack,
      read_data => noblock_obuf_1_2_pipe_read_data,
      write_req => noblock_obuf_1_2_pipe_write_req,
      write_ack => noblock_obuf_1_2_pipe_write_ack,
      write_data => noblock_obuf_1_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_1_3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_1_3",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_1_3_pipe_read_req,
      read_ack => noblock_obuf_1_3_pipe_read_ack,
      read_data => noblock_obuf_1_3_pipe_read_data,
      write_req => noblock_obuf_1_3_pipe_write_req,
      write_ack => noblock_obuf_1_3_pipe_write_ack,
      write_data => noblock_obuf_1_3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_1_4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_1_4",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_1_4_pipe_read_req,
      read_ack => noblock_obuf_1_4_pipe_read_ack,
      read_data => noblock_obuf_1_4_pipe_read_data,
      write_req => noblock_obuf_1_4_pipe_write_req,
      write_ack => noblock_obuf_1_4_pipe_write_ack,
      write_data => noblock_obuf_1_4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_2_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_2_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_2_1_pipe_read_req,
      read_ack => noblock_obuf_2_1_pipe_read_ack,
      read_data => noblock_obuf_2_1_pipe_read_data,
      write_req => noblock_obuf_2_1_pipe_write_req,
      write_ack => noblock_obuf_2_1_pipe_write_ack,
      write_data => noblock_obuf_2_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_2_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_2_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_2_2_pipe_read_req,
      read_ack => noblock_obuf_2_2_pipe_read_ack,
      read_data => noblock_obuf_2_2_pipe_read_data,
      write_req => noblock_obuf_2_2_pipe_write_req,
      write_ack => noblock_obuf_2_2_pipe_write_ack,
      write_data => noblock_obuf_2_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_2_3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_2_3",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_2_3_pipe_read_req,
      read_ack => noblock_obuf_2_3_pipe_read_ack,
      read_data => noblock_obuf_2_3_pipe_read_data,
      write_req => noblock_obuf_2_3_pipe_write_req,
      write_ack => noblock_obuf_2_3_pipe_write_ack,
      write_data => noblock_obuf_2_3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_2_4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_2_4",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_2_4_pipe_read_req,
      read_ack => noblock_obuf_2_4_pipe_read_ack,
      read_data => noblock_obuf_2_4_pipe_read_data,
      write_req => noblock_obuf_2_4_pipe_write_req,
      write_ack => noblock_obuf_2_4_pipe_write_ack,
      write_data => noblock_obuf_2_4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_3_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_3_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_3_1_pipe_read_req,
      read_ack => noblock_obuf_3_1_pipe_read_ack,
      read_data => noblock_obuf_3_1_pipe_read_data,
      write_req => noblock_obuf_3_1_pipe_write_req,
      write_ack => noblock_obuf_3_1_pipe_write_ack,
      write_data => noblock_obuf_3_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_3_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_3_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_3_2_pipe_read_req,
      read_ack => noblock_obuf_3_2_pipe_read_ack,
      read_data => noblock_obuf_3_2_pipe_read_data,
      write_req => noblock_obuf_3_2_pipe_write_req,
      write_ack => noblock_obuf_3_2_pipe_write_ack,
      write_data => noblock_obuf_3_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_3_3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_3_3",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_3_3_pipe_read_req,
      read_ack => noblock_obuf_3_3_pipe_read_ack,
      read_data => noblock_obuf_3_3_pipe_read_data,
      write_req => noblock_obuf_3_3_pipe_write_req,
      write_ack => noblock_obuf_3_3_pipe_write_ack,
      write_data => noblock_obuf_3_3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_3_4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_3_4",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_3_4_pipe_read_req,
      read_ack => noblock_obuf_3_4_pipe_read_ack,
      read_data => noblock_obuf_3_4_pipe_read_data,
      write_req => noblock_obuf_3_4_pipe_write_req,
      write_ack => noblock_obuf_3_4_pipe_write_ack,
      write_data => noblock_obuf_3_4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_4_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_4_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_4_1_pipe_read_req,
      read_ack => noblock_obuf_4_1_pipe_read_ack,
      read_data => noblock_obuf_4_1_pipe_read_data,
      write_req => noblock_obuf_4_1_pipe_write_req,
      write_ack => noblock_obuf_4_1_pipe_write_ack,
      write_data => noblock_obuf_4_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_4_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_4_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_4_2_pipe_read_req,
      read_ack => noblock_obuf_4_2_pipe_read_ack,
      read_data => noblock_obuf_4_2_pipe_read_data,
      write_req => noblock_obuf_4_2_pipe_write_req,
      write_ack => noblock_obuf_4_2_pipe_write_ack,
      write_data => noblock_obuf_4_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_4_3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_4_3",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_4_3_pipe_read_req,
      read_ack => noblock_obuf_4_3_pipe_read_ack,
      read_data => noblock_obuf_4_3_pipe_read_data,
      write_req => noblock_obuf_4_3_pipe_write_req,
      write_ack => noblock_obuf_4_3_pipe_write_ack,
      write_data => noblock_obuf_4_3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  noblock_obuf_4_4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe noblock_obuf_4_4",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 256 --
    )
    port map( -- 
      read_req => noblock_obuf_4_4_pipe_read_req,
      read_ack => noblock_obuf_4_4_pipe_read_ack,
      read_data => noblock_obuf_4_4_pipe_read_data,
      write_req => noblock_obuf_4_4_pipe_write_req,
      write_ack => noblock_obuf_4_4_pipe_write_ack,
      write_data => noblock_obuf_4_4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe out_data_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => out_data_1_pipe_read_req,
      read_ack => out_data_1_pipe_read_ack,
      read_data => out_data_1_pipe_read_data,
      write_req => out_data_1_pipe_write_req,
      write_ack => out_data_1_pipe_write_ack,
      write_data => out_data_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe out_data_2",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => out_data_2_pipe_read_req,
      read_ack => out_data_2_pipe_read_ack,
      read_data => out_data_2_pipe_read_data,
      write_req => out_data_2_pipe_write_req,
      write_ack => out_data_2_pipe_write_ack,
      write_data => out_data_2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe out_data_3",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => out_data_3_pipe_read_req,
      read_ack => out_data_3_pipe_read_ack,
      read_data => out_data_3_pipe_read_data,
      write_req => out_data_3_pipe_write_req,
      write_ack => out_data_3_pipe_write_ack,
      write_data => out_data_3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe out_data_4",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => out_data_4_pipe_read_req,
      read_ack => out_data_4_pipe_read_ack,
      read_data => out_data_4_pipe_read_data,
      write_req => out_data_4_pipe_write_req,
      write_ack => out_data_4_pipe_write_ack,
      write_data => out_data_4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- 
end ahir_system_arch;
